`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09.04.2019 15:57:43
// Design Name: 
// Module Name: top_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: 
// 
//////////////////////////////////////////////////////////////////////////////////

`include "C:\Users\itzka\OneDrive\Documents\Vivado\projects\MNIST_NUMBER_RECOGNITION\src\fpga\rtl\include.v"

`define MaxTestSamples 100

module top_sim(
    );
    
    reg reset;
    reg clock;
    reg [`dataWidth-1:0] in;
    reg in_valid;
    reg [`dataWidth-1:0] in_mem [784:0];
    reg s_axi_awvalid;
    reg [31:0] s_axi_awaddr;
    wire s_axi_awready;
    reg [31:0] s_axi_wdata;
    reg s_axi_wvalid;
    wire s_axi_wready;
    wire s_axi_bvalid;
    reg s_axi_bready;
    wire intr;
    reg [31:0] axiRdData;
    reg [31:0] s_axi_araddr;
    wire [31:0] s_axi_rdata;
    reg s_axi_arvalid;
    wire s_axi_arready;
    wire s_axi_rvalid;
    reg s_axi_rready;
    reg [`dataWidth-1:0] expected;

    wire [31:0] numNeurons[31:1];
    wire [31:0] numWeights[31:1];
    
    assign numNeurons[1] = 30;
    assign numNeurons[2] = 30;
    assign numNeurons[3] = 10;
    assign numNeurons[4] = 10;
    
    assign numWeights[1] = 784;
    assign numWeights[2] = 30;
    assign numWeights[3] = 30;
    assign numWeights[4] = 10;
    
    integer right=0;
    integer wrong=0;
    
    zyNet dut(
    .s_axi_aclk(clock),
    .s_axi_aresetn(reset),
    .s_axi_awaddr(s_axi_awaddr),
    .s_axi_awprot(0),
    .s_axi_awvalid(s_axi_awvalid),
    .s_axi_awready(s_axi_awready),
    .s_axi_wdata(s_axi_wdata),
    .s_axi_wstrb(4'hF),
    .s_axi_wvalid(s_axi_wvalid),
    .s_axi_wready(s_axi_wready),
    .s_axi_bresp(),
    .s_axi_bvalid(s_axi_bvalid),
    .s_axi_bready(s_axi_bready),
    .s_axi_araddr(s_axi_araddr),
    .s_axi_arprot(0),
    .s_axi_arvalid(s_axi_arvalid),
    .s_axi_arready(s_axi_arready),
    .s_axi_rdata(s_axi_rdata),
    .s_axi_rresp(),
    .s_axi_rvalid(s_axi_rvalid),
    .s_axi_rready(s_axi_rready),
    .axis_in_data(in),
    .axis_in_data_valid(in_valid),
    .axis_in_data_ready(),
    .intr(intr)
    );
    
    initial
    begin
        clock = 1'b0;
        s_axi_awvalid = 1'b0;
        s_axi_bready = 1'b0;
        s_axi_wvalid = 1'b0;
        s_axi_arvalid = 1'b0;
    end
        
    always
        #5 clock = ~clock;
    
    always @(posedge clock)
    begin
        s_axi_bready <= s_axi_bvalid;
        s_axi_rready <= s_axi_rvalid;
    end
    
    task writeAxi(
    input [31:0] address,
    input [31:0] data
    );
    begin
        @(posedge clock);
        s_axi_awvalid <= 1'b1;
        s_axi_awaddr <= address;
        s_axi_wdata <= data;
        s_axi_wvalid <= 1'b1;
        wait(s_axi_wready);
        @(posedge clock);
        s_axi_awvalid <= 1'b0;
        s_axi_wvalid <= 1'b0;
        @(posedge clock);
    end
    endtask
    
    task readAxi(
    input [31:0] address
    );
    begin
        @(posedge clock);
        s_axi_arvalid <= 1'b1;
        s_axi_araddr <= address;
        wait(s_axi_arready);
        @(posedge clock);
        s_axi_arvalid <= 1'b0;
        wait(s_axi_rvalid);
        @(posedge clock);
        axiRdData <= s_axi_rdata;
        @(posedge clock);
    end
    endtask
    
    // Define weight file names
    reg [8*20-1:0] weight_files [0:79];
    initial begin
        weight_files[0]  = "w_1_0.mif";  weight_files[1]  = "w_1_1.mif";  weight_files[2]  = "w_1_2.mif";  weight_files[3]  = "w_1_3.mif";
        weight_files[4]  = "w_1_4.mif";  weight_files[5]  = "w_1_5.mif";  weight_files[6]  = "w_1_6.mif";  weight_files[7]  = "w_1_7.mif";
        weight_files[8]  = "w_1_8.mif";  weight_files[9]  = "w_1_9.mif";  weight_files[10] = "w_1_10.mif"; weight_files[11] = "w_1_11.mif";
        weight_files[12] = "w_1_12.mif"; weight_files[13] = "w_1_13.mif"; weight_files[14] = "w_1_14.mif"; weight_files[15] = "w_1_15.mif";
        weight_files[16] = "w_1_16.mif"; weight_files[17] = "w_1_17.mif"; weight_files[18] = "w_1_18.mif"; weight_files[19] = "w_1_19.mif";
        weight_files[20] = "w_1_20.mif"; weight_files[21] = "w_1_21.mif"; weight_files[22] = "w_1_22.mif"; weight_files[23] = "w_1_23.mif";
        weight_files[24] = "w_1_24.mif"; weight_files[25] = "w_1_25.mif"; weight_files[26] = "w_1_26.mif"; weight_files[27] = "w_1_27.mif";
        weight_files[28] = "w_1_28.mif"; weight_files[29] = "w_1_29.mif";
        weight_files[30] = "w_2_0.mif";  weight_files[31] = "w_2_1.mif";  weight_files[32] = "w_2_2.mif";  weight_files[33] = "w_2_3.mif";
        weight_files[34] = "w_2_4.mif";  weight_files[35] = "w_2_5.mif";  weight_files[36] = "w_2_6.mif";  weight_files[37] = "w_2_7.mif";
        weight_files[38] = "w_2_8.mif";  weight_files[39] = "w_2_9.mif";  weight_files[40] = "w_2_10.mif"; weight_files[41] = "w_2_11.mif";
        weight_files[42] = "w_2_12.mif"; weight_files[43] = "w_2_13.mif"; weight_files[44] = "w_2_14.mif"; weight_files[45] = "w_2_15.mif";
        weight_files[46] = "w_2_16.mif"; weight_files[47] = "w_2_17.mif"; weight_files[48] = "w_2_18.mif"; weight_files[49] = "w_2_19.mif";
        weight_files[50] = "w_2_20.mif"; weight_files[51] = "w_2_21.mif"; weight_files[52] = "w_2_22.mif"; weight_files[53] = "w_2_23.mif";
        weight_files[54] = "w_2_24.mif"; weight_files[55] = "w_2_25.mif"; weight_files[56] = "w_2_26.mif"; weight_files[57] = "w_2_27.mif";
        weight_files[58] = "w_2_28.mif"; weight_files[59] = "w_2_29.mif";
        weight_files[60] = "w_3_0.mif";  weight_files[61] = "w_3_1.mif";  weight_files[62] = "w_3_2.mif";  weight_files[63] = "w_3_3.mif";
        weight_files[64] = "w_3_4.mif";  weight_files[65] = "w_3_5.mif";  weight_files[66] = "w_3_6.mif";  weight_files[67] = "w_3_7.mif";
        weight_files[68] = "w_3_8.mif";  weight_files[69] = "w_3_9.mif";
        weight_files[70] = "w_4_0.mif";  weight_files[71] = "w_4_1.mif";  weight_files[72] = "w_4_2.mif";  weight_files[73] = "w_4_3.mif";
        weight_files[74] = "w_4_4.mif";  weight_files[75] = "w_4_5.mif";  weight_files[76] = "w_4_6.mif";  weight_files[77] = "w_4_7.mif";
        weight_files[78] = "w_4_8.mif";  weight_files[79] = "w_4_9.mif";
    end

    // Define bias file names
    reg [8*20-1:0] bias_files [0:79];
    initial begin
        bias_files[0]  = "b_1_0.mif";  bias_files[1]  = "b_1_1.mif";  bias_files[2]  = "b_1_2.mif";  bias_files[3]  = "b_1_3.mif";
        bias_files[4]  = "b_1_4.mif";  bias_files[5]  = "b_1_5.mif";  bias_files[6]  = "b_1_6.mif";  bias_files[7]  = "b_1_7.mif";
        bias_files[8]  = "b_1_8.mif";  bias_files[9]  = "b_1_9.mif";  bias_files[10] = "b_1_10.mif"; bias_files[11] = "b_1_11.mif";
        bias_files[12] = "b_1_12.mif"; bias_files[13] = "b_1_13.mif"; bias_files[14] = "b_1_14.mif"; bias_files[15] = "b_1_15.mif";
        bias_files[16] = "b_1_16.mif"; bias_files[17] = "b_1_17.mif"; bias_files[18] = "b_1_18.mif"; bias_files[19] = "b_1_19.mif";
        bias_files[20] = "b_1_20.mif"; bias_files[21] = "b_1_21.mif"; bias_files[22] = "b_1_22.mif"; bias_files[23] = "b_1_23.mif";
        bias_files[24] = "b_1_24.mif"; bias_files[25] = "b_1_25.mif"; bias_files[26] = "b_1_26.mif"; bias_files[27] = "b_1_27.mif";
        bias_files[28] = "b_1_28.mif"; bias_files[29] = "b_1_29.mif";
        bias_files[30] = "b_2_0.mif";  bias_files[31] = "b_2_1.mif";  bias_files[32] = "b_2_2.mif";  bias_files[33] = "b_2_3.mif";
        bias_files[34] = "b_2_4.mif";  bias_files[35] = "b_2_5.mif";  bias_files[36] = "b_2_6.mif";  bias_files[37] = "b_2_7.mif";
        bias_files[38] = "b_2_8.mif";  bias_files[39] = "b_2_9.mif";  bias_files[40] = "b_2_10.mif"; bias_files[41] = "b_2_11.mif";
        bias_files[42] = "b_2_12.mif"; bias_files[43] = "b_2_13.mif"; bias_files[44] = "b_2_14.mif"; bias_files[45] = "b_2_15.mif";
        bias_files[46] = "b_2_16.mif"; bias_files[47] = "b_2_17.mif"; bias_files[48] = "b_2_18.mif"; bias_files[49] = "b_2_19.mif";
        bias_files[50] = "b_2_20.mif"; bias_files[51] = "b_2_21.mif"; bias_files[52] = "b_2_22.mif"; bias_files[53] = "b_2_23.mif";
        bias_files[54] = "b_2_24.mif"; bias_files[55] = "b_2_25.mif"; bias_files[56] = "b_2_26.mif"; bias_files[57] = "b_2_27.mif";
        bias_files[58] = "b_2_28.mif"; bias_files[59] = "b_2_29.mif";
        bias_files[60] = "b_3_0.mif";  bias_files[61] = "b_3_1.mif";  bias_files[62] = "b_3_2.mif";  bias_files[63] = "b_3_3.mif";
        bias_files[64] = "b_3_4.mif";  bias_files[65] = "b_3_5.mif";  bias_files[66] = "b_3_6.mif";  bias_files[67] = "b_3_7.mif";
        bias_files[68] = "b_3_8.mif";  bias_files[69] = "b_3_9.mif";
        bias_files[70] = "b_4_0.mif";  bias_files[71] = "b_4_1.mif";  bias_files[72] = "b_4_2.mif";  bias_files[73] = "b_4_3.mif";
        bias_files[74] = "b_4_4.mif";  bias_files[75] = "b_4_5.mif";  bias_files[76] = "b_4_6.mif";  bias_files[77] = "b_4_7.mif";
        bias_files[78] = "b_4_8.mif";  bias_files[79] = "b_4_9.mif";
    end

    task configWeights();
    integer j, k, t;
    integer file_idx;
    reg [`dataWidth:0] config_mem [783:0];
    begin
        @(posedge clock);
        file_idx = 0;
        for(k=1; k<=`numLayers; k=k+1)
        begin
            writeAxi(12, k); // Write layer number
            for(j=0; j<numNeurons[k]; j=j+1)
            begin
                $readmemb(weight_files[file_idx], config_mem);
                writeAxi(16, j); // Write neuron number
                for (t=0; t<numWeights[k]; t=t+1) begin
                    writeAxi(0, {15'd0, config_mem[t]});
                end
                file_idx = file_idx + 1;
            end
        end
    end
    endtask
    
    task configBias();
    integer j, k;
    integer file_idx;
    reg [31:0] bias[0:0];
    begin
        @(posedge clock);
        file_idx = 0;
        for(k=1; k<=`numLayers; k=k+1)
        begin
            writeAxi(12, k); // Write layer number
            for(j=0; j<numNeurons[k]; j=j+1)
            begin
                $readmemb(bias_files[file_idx], bias);
                writeAxi(16, j); // Write neuron number
                writeAxi(4, {15'd0, bias[0]});
                file_idx = file_idx + 1;
            end
        end
    end
    endtask
    
    // Define test data file names
    reg [8*20-1:0] test_data_files [0:9999];
    initial begin
        test_data_files[0] = "test_data_0000.txt";
test_data_files[1] = "test_data_0001.txt";
test_data_files[2] = "test_data_0002.txt";
test_data_files[3] = "test_data_0003.txt";
test_data_files[4] = "test_data_0004.txt";
test_data_files[5] = "test_data_0005.txt";
test_data_files[6] = "test_data_0006.txt";
test_data_files[7] = "test_data_0007.txt";
test_data_files[8] = "test_data_0008.txt";
test_data_files[9] = "test_data_0009.txt";
test_data_files[10] = "test_data_0010.txt";
test_data_files[11] = "test_data_0011.txt";
test_data_files[12] = "test_data_0012.txt";
test_data_files[13] = "test_data_0013.txt";
test_data_files[14] = "test_data_0014.txt";
test_data_files[15] = "test_data_0015.txt";
test_data_files[16] = "test_data_0016.txt";
test_data_files[17] = "test_data_0017.txt";
test_data_files[18] = "test_data_0018.txt";
test_data_files[19] = "test_data_0019.txt";
test_data_files[20] = "test_data_0020.txt";
test_data_files[21] = "test_data_0021.txt";
test_data_files[22] = "test_data_0022.txt";
test_data_files[23] = "test_data_0023.txt";
test_data_files[24] = "test_data_0024.txt";
test_data_files[25] = "test_data_0025.txt";
test_data_files[26] = "test_data_0026.txt";
test_data_files[27] = "test_data_0027.txt";
test_data_files[28] = "test_data_0028.txt";
test_data_files[29] = "test_data_0029.txt";
test_data_files[30] = "test_data_0030.txt";
test_data_files[31] = "test_data_0031.txt";
test_data_files[32] = "test_data_0032.txt";
test_data_files[33] = "test_data_0033.txt";
test_data_files[34] = "test_data_0034.txt";
test_data_files[35] = "test_data_0035.txt";
test_data_files[36] = "test_data_0036.txt";
test_data_files[37] = "test_data_0037.txt";
test_data_files[38] = "test_data_0038.txt";
test_data_files[39] = "test_data_0039.txt";
test_data_files[40] = "test_data_0040.txt";
test_data_files[41] = "test_data_0041.txt";
test_data_files[42] = "test_data_0042.txt";
test_data_files[43] = "test_data_0043.txt";
test_data_files[44] = "test_data_0044.txt";
test_data_files[45] = "test_data_0045.txt";
test_data_files[46] = "test_data_0046.txt";
test_data_files[47] = "test_data_0047.txt";
test_data_files[48] = "test_data_0048.txt";
test_data_files[49] = "test_data_0049.txt";
test_data_files[50] = "test_data_0050.txt";
test_data_files[51] = "test_data_0051.txt";
test_data_files[52] = "test_data_0052.txt";
test_data_files[53] = "test_data_0053.txt";
test_data_files[54] = "test_data_0054.txt";
test_data_files[55] = "test_data_0055.txt";
test_data_files[56] = "test_data_0056.txt";
test_data_files[57] = "test_data_0057.txt";
test_data_files[58] = "test_data_0058.txt";
test_data_files[59] = "test_data_0059.txt";
test_data_files[60] = "test_data_0060.txt";
test_data_files[61] = "test_data_0061.txt";
test_data_files[62] = "test_data_0062.txt";
test_data_files[63] = "test_data_0063.txt";
test_data_files[64] = "test_data_0064.txt";
test_data_files[65] = "test_data_0065.txt";
test_data_files[66] = "test_data_0066.txt";
test_data_files[67] = "test_data_0067.txt";
test_data_files[68] = "test_data_0068.txt";
test_data_files[69] = "test_data_0069.txt";
test_data_files[70] = "test_data_0070.txt";
test_data_files[71] = "test_data_0071.txt";
test_data_files[72] = "test_data_0072.txt";
test_data_files[73] = "test_data_0073.txt";
test_data_files[74] = "test_data_0074.txt";
test_data_files[75] = "test_data_0075.txt";
test_data_files[76] = "test_data_0076.txt";
test_data_files[77] = "test_data_0077.txt";
test_data_files[78] = "test_data_0078.txt";
test_data_files[79] = "test_data_0079.txt";
test_data_files[80] = "test_data_0080.txt";
test_data_files[81] = "test_data_0081.txt";
test_data_files[82] = "test_data_0082.txt";
test_data_files[83] = "test_data_0083.txt";
test_data_files[84] = "test_data_0084.txt";
test_data_files[85] = "test_data_0085.txt";
test_data_files[86] = "test_data_0086.txt";
test_data_files[87] = "test_data_0087.txt";
test_data_files[88] = "test_data_0088.txt";
test_data_files[89] = "test_data_0089.txt";
test_data_files[90] = "test_data_0090.txt";
test_data_files[91] = "test_data_0091.txt";
test_data_files[92] = "test_data_0092.txt";
test_data_files[93] = "test_data_0093.txt";
test_data_files[94] = "test_data_0094.txt";
test_data_files[95] = "test_data_0095.txt";
test_data_files[96] = "test_data_0096.txt";
test_data_files[97] = "test_data_0097.txt";
test_data_files[98] = "test_data_0098.txt";
test_data_files[99] = "test_data_0099.txt";
test_data_files[100] = "test_data_0100.txt";
test_data_files[101] = "test_data_0101.txt";
test_data_files[102] = "test_data_0102.txt";
test_data_files[103] = "test_data_0103.txt";
test_data_files[104] = "test_data_0104.txt";
test_data_files[105] = "test_data_0105.txt";
test_data_files[106] = "test_data_0106.txt";
test_data_files[107] = "test_data_0107.txt";
test_data_files[108] = "test_data_0108.txt";
test_data_files[109] = "test_data_0109.txt";
test_data_files[110] = "test_data_0110.txt";
test_data_files[111] = "test_data_0111.txt";
test_data_files[112] = "test_data_0112.txt";
test_data_files[113] = "test_data_0113.txt";
test_data_files[114] = "test_data_0114.txt";
test_data_files[115] = "test_data_0115.txt";
test_data_files[116] = "test_data_0116.txt";
test_data_files[117] = "test_data_0117.txt";
test_data_files[118] = "test_data_0118.txt";
test_data_files[119] = "test_data_0119.txt";
test_data_files[120] = "test_data_0120.txt";
test_data_files[121] = "test_data_0121.txt";
test_data_files[122] = "test_data_0122.txt";
test_data_files[123] = "test_data_0123.txt";
test_data_files[124] = "test_data_0124.txt";
test_data_files[125] = "test_data_0125.txt";
test_data_files[126] = "test_data_0126.txt";
test_data_files[127] = "test_data_0127.txt";
test_data_files[128] = "test_data_0128.txt";
test_data_files[129] = "test_data_0129.txt";
test_data_files[130] = "test_data_0130.txt";
test_data_files[131] = "test_data_0131.txt";
test_data_files[132] = "test_data_0132.txt";
test_data_files[133] = "test_data_0133.txt";
test_data_files[134] = "test_data_0134.txt";
test_data_files[135] = "test_data_0135.txt";
test_data_files[136] = "test_data_0136.txt";
test_data_files[137] = "test_data_0137.txt";
test_data_files[138] = "test_data_0138.txt";
test_data_files[139] = "test_data_0139.txt";
test_data_files[140] = "test_data_0140.txt";
test_data_files[141] = "test_data_0141.txt";
test_data_files[142] = "test_data_0142.txt";
test_data_files[143] = "test_data_0143.txt";
test_data_files[144] = "test_data_0144.txt";
test_data_files[145] = "test_data_0145.txt";
test_data_files[146] = "test_data_0146.txt";
test_data_files[147] = "test_data_0147.txt";
test_data_files[148] = "test_data_0148.txt";
test_data_files[149] = "test_data_0149.txt";
test_data_files[150] = "test_data_0150.txt";
test_data_files[151] = "test_data_0151.txt";
test_data_files[152] = "test_data_0152.txt";
test_data_files[153] = "test_data_0153.txt";
test_data_files[154] = "test_data_0154.txt";
test_data_files[155] = "test_data_0155.txt";
test_data_files[156] = "test_data_0156.txt";
test_data_files[157] = "test_data_0157.txt";
test_data_files[158] = "test_data_0158.txt";
test_data_files[159] = "test_data_0159.txt";
test_data_files[160] = "test_data_0160.txt";
test_data_files[161] = "test_data_0161.txt";
test_data_files[162] = "test_data_0162.txt";
test_data_files[163] = "test_data_0163.txt";
test_data_files[164] = "test_data_0164.txt";
test_data_files[165] = "test_data_0165.txt";
test_data_files[166] = "test_data_0166.txt";
test_data_files[167] = "test_data_0167.txt";
test_data_files[168] = "test_data_0168.txt";
test_data_files[169] = "test_data_0169.txt";
test_data_files[170] = "test_data_0170.txt";
test_data_files[171] = "test_data_0171.txt";
test_data_files[172] = "test_data_0172.txt";
test_data_files[173] = "test_data_0173.txt";
test_data_files[174] = "test_data_0174.txt";
test_data_files[175] = "test_data_0175.txt";
test_data_files[176] = "test_data_0176.txt";
test_data_files[177] = "test_data_0177.txt";
test_data_files[178] = "test_data_0178.txt";
test_data_files[179] = "test_data_0179.txt";
test_data_files[180] = "test_data_0180.txt";
test_data_files[181] = "test_data_0181.txt";
test_data_files[182] = "test_data_0182.txt";
test_data_files[183] = "test_data_0183.txt";
test_data_files[184] = "test_data_0184.txt";
test_data_files[185] = "test_data_0185.txt";
test_data_files[186] = "test_data_0186.txt";
test_data_files[187] = "test_data_0187.txt";
test_data_files[188] = "test_data_0188.txt";
test_data_files[189] = "test_data_0189.txt";
test_data_files[190] = "test_data_0190.txt";
test_data_files[191] = "test_data_0191.txt";
test_data_files[192] = "test_data_0192.txt";
test_data_files[193] = "test_data_0193.txt";
test_data_files[194] = "test_data_0194.txt";
test_data_files[195] = "test_data_0195.txt";
test_data_files[196] = "test_data_0196.txt";
test_data_files[197] = "test_data_0197.txt";
test_data_files[198] = "test_data_0198.txt";
test_data_files[199] = "test_data_0199.txt";
test_data_files[200] = "test_data_0200.txt";
test_data_files[201] = "test_data_0201.txt";
test_data_files[202] = "test_data_0202.txt";
test_data_files[203] = "test_data_0203.txt";
test_data_files[204] = "test_data_0204.txt";
test_data_files[205] = "test_data_0205.txt";
test_data_files[206] = "test_data_0206.txt";
test_data_files[207] = "test_data_0207.txt";
test_data_files[208] = "test_data_0208.txt";
test_data_files[209] = "test_data_0209.txt";
test_data_files[210] = "test_data_0210.txt";
test_data_files[211] = "test_data_0211.txt";
test_data_files[212] = "test_data_0212.txt";
test_data_files[213] = "test_data_0213.txt";
test_data_files[214] = "test_data_0214.txt";
test_data_files[215] = "test_data_0215.txt";
test_data_files[216] = "test_data_0216.txt";
test_data_files[217] = "test_data_0217.txt";
test_data_files[218] = "test_data_0218.txt";
test_data_files[219] = "test_data_0219.txt";
test_data_files[220] = "test_data_0220.txt";
test_data_files[221] = "test_data_0221.txt";
test_data_files[222] = "test_data_0222.txt";
test_data_files[223] = "test_data_0223.txt";
test_data_files[224] = "test_data_0224.txt";
test_data_files[225] = "test_data_0225.txt";
test_data_files[226] = "test_data_0226.txt";
test_data_files[227] = "test_data_0227.txt";
test_data_files[228] = "test_data_0228.txt";
test_data_files[229] = "test_data_0229.txt";
test_data_files[230] = "test_data_0230.txt";
test_data_files[231] = "test_data_0231.txt";
test_data_files[232] = "test_data_0232.txt";
test_data_files[233] = "test_data_0233.txt";
test_data_files[234] = "test_data_0234.txt";
test_data_files[235] = "test_data_0235.txt";
test_data_files[236] = "test_data_0236.txt";
test_data_files[237] = "test_data_0237.txt";
test_data_files[238] = "test_data_0238.txt";
test_data_files[239] = "test_data_0239.txt";
test_data_files[240] = "test_data_0240.txt";
test_data_files[241] = "test_data_0241.txt";
test_data_files[242] = "test_data_0242.txt";
test_data_files[243] = "test_data_0243.txt";
test_data_files[244] = "test_data_0244.txt";
test_data_files[245] = "test_data_0245.txt";
test_data_files[246] = "test_data_0246.txt";
test_data_files[247] = "test_data_0247.txt";
test_data_files[248] = "test_data_0248.txt";
test_data_files[249] = "test_data_0249.txt";
test_data_files[250] = "test_data_0250.txt";
test_data_files[251] = "test_data_0251.txt";
test_data_files[252] = "test_data_0252.txt";
test_data_files[253] = "test_data_0253.txt";
test_data_files[254] = "test_data_0254.txt";
test_data_files[255] = "test_data_0255.txt";
test_data_files[256] = "test_data_0256.txt";
test_data_files[257] = "test_data_0257.txt";
test_data_files[258] = "test_data_0258.txt";
test_data_files[259] = "test_data_0259.txt";
test_data_files[260] = "test_data_0260.txt";
test_data_files[261] = "test_data_0261.txt";
test_data_files[262] = "test_data_0262.txt";
test_data_files[263] = "test_data_0263.txt";
test_data_files[264] = "test_data_0264.txt";
test_data_files[265] = "test_data_0265.txt";
test_data_files[266] = "test_data_0266.txt";
test_data_files[267] = "test_data_0267.txt";
test_data_files[268] = "test_data_0268.txt";
test_data_files[269] = "test_data_0269.txt";
test_data_files[270] = "test_data_0270.txt";
test_data_files[271] = "test_data_0271.txt";
test_data_files[272] = "test_data_0272.txt";
test_data_files[273] = "test_data_0273.txt";
test_data_files[274] = "test_data_0274.txt";
test_data_files[275] = "test_data_0275.txt";
test_data_files[276] = "test_data_0276.txt";
test_data_files[277] = "test_data_0277.txt";
test_data_files[278] = "test_data_0278.txt";
test_data_files[279] = "test_data_0279.txt";
test_data_files[280] = "test_data_0280.txt";
test_data_files[281] = "test_data_0281.txt";
test_data_files[282] = "test_data_0282.txt";
test_data_files[283] = "test_data_0283.txt";
test_data_files[284] = "test_data_0284.txt";
test_data_files[285] = "test_data_0285.txt";
test_data_files[286] = "test_data_0286.txt";
test_data_files[287] = "test_data_0287.txt";
test_data_files[288] = "test_data_0288.txt";
test_data_files[289] = "test_data_0289.txt";
test_data_files[290] = "test_data_0290.txt";
test_data_files[291] = "test_data_0291.txt";
test_data_files[292] = "test_data_0292.txt";
test_data_files[293] = "test_data_0293.txt";
test_data_files[294] = "test_data_0294.txt";
test_data_files[295] = "test_data_0295.txt";
test_data_files[296] = "test_data_0296.txt";
test_data_files[297] = "test_data_0297.txt";
test_data_files[298] = "test_data_0298.txt";
test_data_files[299] = "test_data_0299.txt";
test_data_files[300] = "test_data_0300.txt";
test_data_files[301] = "test_data_0301.txt";
test_data_files[302] = "test_data_0302.txt";
test_data_files[303] = "test_data_0303.txt";
test_data_files[304] = "test_data_0304.txt";
test_data_files[305] = "test_data_0305.txt";
test_data_files[306] = "test_data_0306.txt";
test_data_files[307] = "test_data_0307.txt";
test_data_files[308] = "test_data_0308.txt";
test_data_files[309] = "test_data_0309.txt";
test_data_files[310] = "test_data_0310.txt";
test_data_files[311] = "test_data_0311.txt";
test_data_files[312] = "test_data_0312.txt";
test_data_files[313] = "test_data_0313.txt";
test_data_files[314] = "test_data_0314.txt";
test_data_files[315] = "test_data_0315.txt";
test_data_files[316] = "test_data_0316.txt";
test_data_files[317] = "test_data_0317.txt";
test_data_files[318] = "test_data_0318.txt";
test_data_files[319] = "test_data_0319.txt";
test_data_files[320] = "test_data_0320.txt";
test_data_files[321] = "test_data_0321.txt";
test_data_files[322] = "test_data_0322.txt";
test_data_files[323] = "test_data_0323.txt";
test_data_files[324] = "test_data_0324.txt";
test_data_files[325] = "test_data_0325.txt";
test_data_files[326] = "test_data_0326.txt";
test_data_files[327] = "test_data_0327.txt";
test_data_files[328] = "test_data_0328.txt";
test_data_files[329] = "test_data_0329.txt";
test_data_files[330] = "test_data_0330.txt";
test_data_files[331] = "test_data_0331.txt";
test_data_files[332] = "test_data_0332.txt";
test_data_files[333] = "test_data_0333.txt";
test_data_files[334] = "test_data_0334.txt";
test_data_files[335] = "test_data_0335.txt";
test_data_files[336] = "test_data_0336.txt";
test_data_files[337] = "test_data_0337.txt";
test_data_files[338] = "test_data_0338.txt";
test_data_files[339] = "test_data_0339.txt";
test_data_files[340] = "test_data_0340.txt";
test_data_files[341] = "test_data_0341.txt";
test_data_files[342] = "test_data_0342.txt";
test_data_files[343] = "test_data_0343.txt";
test_data_files[344] = "test_data_0344.txt";
test_data_files[345] = "test_data_0345.txt";
test_data_files[346] = "test_data_0346.txt";
test_data_files[347] = "test_data_0347.txt";
test_data_files[348] = "test_data_0348.txt";
test_data_files[349] = "test_data_0349.txt";
test_data_files[350] = "test_data_0350.txt";
test_data_files[351] = "test_data_0351.txt";
test_data_files[352] = "test_data_0352.txt";
test_data_files[353] = "test_data_0353.txt";
test_data_files[354] = "test_data_0354.txt";
test_data_files[355] = "test_data_0355.txt";
test_data_files[356] = "test_data_0356.txt";
test_data_files[357] = "test_data_0357.txt";
test_data_files[358] = "test_data_0358.txt";
test_data_files[359] = "test_data_0359.txt";
test_data_files[360] = "test_data_0360.txt";
test_data_files[361] = "test_data_0361.txt";
test_data_files[362] = "test_data_0362.txt";
test_data_files[363] = "test_data_0363.txt";
test_data_files[364] = "test_data_0364.txt";
test_data_files[365] = "test_data_0365.txt";
test_data_files[366] = "test_data_0366.txt";
test_data_files[367] = "test_data_0367.txt";
test_data_files[368] = "test_data_0368.txt";
test_data_files[369] = "test_data_0369.txt";
test_data_files[370] = "test_data_0370.txt";
test_data_files[371] = "test_data_0371.txt";
test_data_files[372] = "test_data_0372.txt";
test_data_files[373] = "test_data_0373.txt";
test_data_files[374] = "test_data_0374.txt";
test_data_files[375] = "test_data_0375.txt";
test_data_files[376] = "test_data_0376.txt";
test_data_files[377] = "test_data_0377.txt";
test_data_files[378] = "test_data_0378.txt";
test_data_files[379] = "test_data_0379.txt";
test_data_files[380] = "test_data_0380.txt";
test_data_files[381] = "test_data_0381.txt";
test_data_files[382] = "test_data_0382.txt";
test_data_files[383] = "test_data_0383.txt";
test_data_files[384] = "test_data_0384.txt";
test_data_files[385] = "test_data_0385.txt";
test_data_files[386] = "test_data_0386.txt";
test_data_files[387] = "test_data_0387.txt";
test_data_files[388] = "test_data_0388.txt";
test_data_files[389] = "test_data_0389.txt";
test_data_files[390] = "test_data_0390.txt";
test_data_files[391] = "test_data_0391.txt";
test_data_files[392] = "test_data_0392.txt";
test_data_files[393] = "test_data_0393.txt";
test_data_files[394] = "test_data_0394.txt";
test_data_files[395] = "test_data_0395.txt";
test_data_files[396] = "test_data_0396.txt";
test_data_files[397] = "test_data_0397.txt";
test_data_files[398] = "test_data_0398.txt";
test_data_files[399] = "test_data_0399.txt";
test_data_files[400] = "test_data_0400.txt";
test_data_files[401] = "test_data_0401.txt";
test_data_files[402] = "test_data_0402.txt";
test_data_files[403] = "test_data_0403.txt";
test_data_files[404] = "test_data_0404.txt";
test_data_files[405] = "test_data_0405.txt";
test_data_files[406] = "test_data_0406.txt";
test_data_files[407] = "test_data_0407.txt";
test_data_files[408] = "test_data_0408.txt";
test_data_files[409] = "test_data_0409.txt";
test_data_files[410] = "test_data_0410.txt";
test_data_files[411] = "test_data_0411.txt";
test_data_files[412] = "test_data_0412.txt";
test_data_files[413] = "test_data_0413.txt";
test_data_files[414] = "test_data_0414.txt";
test_data_files[415] = "test_data_0415.txt";
test_data_files[416] = "test_data_0416.txt";
test_data_files[417] = "test_data_0417.txt";
test_data_files[418] = "test_data_0418.txt";
test_data_files[419] = "test_data_0419.txt";
test_data_files[420] = "test_data_0420.txt";
test_data_files[421] = "test_data_0421.txt";
test_data_files[422] = "test_data_0422.txt";
test_data_files[423] = "test_data_0423.txt";
test_data_files[424] = "test_data_0424.txt";
test_data_files[425] = "test_data_0425.txt";
test_data_files[426] = "test_data_0426.txt";
test_data_files[427] = "test_data_0427.txt";
test_data_files[428] = "test_data_0428.txt";
test_data_files[429] = "test_data_0429.txt";
test_data_files[430] = "test_data_0430.txt";
test_data_files[431] = "test_data_0431.txt";
test_data_files[432] = "test_data_0432.txt";
test_data_files[433] = "test_data_0433.txt";
test_data_files[434] = "test_data_0434.txt";
test_data_files[435] = "test_data_0435.txt";
test_data_files[436] = "test_data_0436.txt";
test_data_files[437] = "test_data_0437.txt";
test_data_files[438] = "test_data_0438.txt";
test_data_files[439] = "test_data_0439.txt";
test_data_files[440] = "test_data_0440.txt";
test_data_files[441] = "test_data_0441.txt";
test_data_files[442] = "test_data_0442.txt";
test_data_files[443] = "test_data_0443.txt";
test_data_files[444] = "test_data_0444.txt";
test_data_files[445] = "test_data_0445.txt";
test_data_files[446] = "test_data_0446.txt";
test_data_files[447] = "test_data_0447.txt";
test_data_files[448] = "test_data_0448.txt";
test_data_files[449] = "test_data_0449.txt";
test_data_files[450] = "test_data_0450.txt";
test_data_files[451] = "test_data_0451.txt";
test_data_files[452] = "test_data_0452.txt";
test_data_files[453] = "test_data_0453.txt";
test_data_files[454] = "test_data_0454.txt";
test_data_files[455] = "test_data_0455.txt";
test_data_files[456] = "test_data_0456.txt";
test_data_files[457] = "test_data_0457.txt";
test_data_files[458] = "test_data_0458.txt";
test_data_files[459] = "test_data_0459.txt";
test_data_files[460] = "test_data_0460.txt";
test_data_files[461] = "test_data_0461.txt";
test_data_files[462] = "test_data_0462.txt";
test_data_files[463] = "test_data_0463.txt";
test_data_files[464] = "test_data_0464.txt";
test_data_files[465] = "test_data_0465.txt";
test_data_files[466] = "test_data_0466.txt";
test_data_files[467] = "test_data_0467.txt";
test_data_files[468] = "test_data_0468.txt";
test_data_files[469] = "test_data_0469.txt";
test_data_files[470] = "test_data_0470.txt";
test_data_files[471] = "test_data_0471.txt";
test_data_files[472] = "test_data_0472.txt";
test_data_files[473] = "test_data_0473.txt";
test_data_files[474] = "test_data_0474.txt";
test_data_files[475] = "test_data_0475.txt";
test_data_files[476] = "test_data_0476.txt";
test_data_files[477] = "test_data_0477.txt";
test_data_files[478] = "test_data_0478.txt";
test_data_files[479] = "test_data_0479.txt";
test_data_files[480] = "test_data_0480.txt";
test_data_files[481] = "test_data_0481.txt";
test_data_files[482] = "test_data_0482.txt";
test_data_files[483] = "test_data_0483.txt";
test_data_files[484] = "test_data_0484.txt";
test_data_files[485] = "test_data_0485.txt";
test_data_files[486] = "test_data_0486.txt";
test_data_files[487] = "test_data_0487.txt";
test_data_files[488] = "test_data_0488.txt";
test_data_files[489] = "test_data_0489.txt";
test_data_files[490] = "test_data_0490.txt";
test_data_files[491] = "test_data_0491.txt";
test_data_files[492] = "test_data_0492.txt";
test_data_files[493] = "test_data_0493.txt";
test_data_files[494] = "test_data_0494.txt";
test_data_files[495] = "test_data_0495.txt";
test_data_files[496] = "test_data_0496.txt";
test_data_files[497] = "test_data_0497.txt";
test_data_files[498] = "test_data_0498.txt";
test_data_files[499] = "test_data_0499.txt";
test_data_files[500] = "test_data_0500.txt";
test_data_files[501] = "test_data_0501.txt";
test_data_files[502] = "test_data_0502.txt";
test_data_files[503] = "test_data_0503.txt";
test_data_files[504] = "test_data_0504.txt";
test_data_files[505] = "test_data_0505.txt";
test_data_files[506] = "test_data_0506.txt";
test_data_files[507] = "test_data_0507.txt";
test_data_files[508] = "test_data_0508.txt";
test_data_files[509] = "test_data_0509.txt";
test_data_files[510] = "test_data_0510.txt";
test_data_files[511] = "test_data_0511.txt";
test_data_files[512] = "test_data_0512.txt";
test_data_files[513] = "test_data_0513.txt";
test_data_files[514] = "test_data_0514.txt";
test_data_files[515] = "test_data_0515.txt";
test_data_files[516] = "test_data_0516.txt";
test_data_files[517] = "test_data_0517.txt";
test_data_files[518] = "test_data_0518.txt";
test_data_files[519] = "test_data_0519.txt";
test_data_files[520] = "test_data_0520.txt";
test_data_files[521] = "test_data_0521.txt";
test_data_files[522] = "test_data_0522.txt";
test_data_files[523] = "test_data_0523.txt";
test_data_files[524] = "test_data_0524.txt";
test_data_files[525] = "test_data_0525.txt";
test_data_files[526] = "test_data_0526.txt";
test_data_files[527] = "test_data_0527.txt";
test_data_files[528] = "test_data_0528.txt";
test_data_files[529] = "test_data_0529.txt";
test_data_files[530] = "test_data_0530.txt";
test_data_files[531] = "test_data_0531.txt";
test_data_files[532] = "test_data_0532.txt";
test_data_files[533] = "test_data_0533.txt";
test_data_files[534] = "test_data_0534.txt";
test_data_files[535] = "test_data_0535.txt";
test_data_files[536] = "test_data_0536.txt";
test_data_files[537] = "test_data_0537.txt";
test_data_files[538] = "test_data_0538.txt";
test_data_files[539] = "test_data_0539.txt";
test_data_files[540] = "test_data_0540.txt";
test_data_files[541] = "test_data_0541.txt";
test_data_files[542] = "test_data_0542.txt";
test_data_files[543] = "test_data_0543.txt";
test_data_files[544] = "test_data_0544.txt";
test_data_files[545] = "test_data_0545.txt";
test_data_files[546] = "test_data_0546.txt";
test_data_files[547] = "test_data_0547.txt";
test_data_files[548] = "test_data_0548.txt";
test_data_files[549] = "test_data_0549.txt";
test_data_files[550] = "test_data_0550.txt";
test_data_files[551] = "test_data_0551.txt";
test_data_files[552] = "test_data_0552.txt";
test_data_files[553] = "test_data_0553.txt";
test_data_files[554] = "test_data_0554.txt";
test_data_files[555] = "test_data_0555.txt";
test_data_files[556] = "test_data_0556.txt";
test_data_files[557] = "test_data_0557.txt";
test_data_files[558] = "test_data_0558.txt";
test_data_files[559] = "test_data_0559.txt";
test_data_files[560] = "test_data_0560.txt";
test_data_files[561] = "test_data_0561.txt";
test_data_files[562] = "test_data_0562.txt";
test_data_files[563] = "test_data_0563.txt";
test_data_files[564] = "test_data_0564.txt";
test_data_files[565] = "test_data_0565.txt";
test_data_files[566] = "test_data_0566.txt";
test_data_files[567] = "test_data_0567.txt";
test_data_files[568] = "test_data_0568.txt";
test_data_files[569] = "test_data_0569.txt";
test_data_files[570] = "test_data_0570.txt";
test_data_files[571] = "test_data_0571.txt";
test_data_files[572] = "test_data_0572.txt";
test_data_files[573] = "test_data_0573.txt";
test_data_files[574] = "test_data_0574.txt";
test_data_files[575] = "test_data_0575.txt";
test_data_files[576] = "test_data_0576.txt";
test_data_files[577] = "test_data_0577.txt";
test_data_files[578] = "test_data_0578.txt";
test_data_files[579] = "test_data_0579.txt";
test_data_files[580] = "test_data_0580.txt";
test_data_files[581] = "test_data_0581.txt";
test_data_files[582] = "test_data_0582.txt";
test_data_files[583] = "test_data_0583.txt";
test_data_files[584] = "test_data_0584.txt";
test_data_files[585] = "test_data_0585.txt";
test_data_files[586] = "test_data_0586.txt";
test_data_files[587] = "test_data_0587.txt";
test_data_files[588] = "test_data_0588.txt";
test_data_files[589] = "test_data_0589.txt";
test_data_files[590] = "test_data_0590.txt";
test_data_files[591] = "test_data_0591.txt";
test_data_files[592] = "test_data_0592.txt";
test_data_files[593] = "test_data_0593.txt";
test_data_files[594] = "test_data_0594.txt";
test_data_files[595] = "test_data_0595.txt";
test_data_files[596] = "test_data_0596.txt";
test_data_files[597] = "test_data_0597.txt";
test_data_files[598] = "test_data_0598.txt";
test_data_files[599] = "test_data_0599.txt";
test_data_files[600] = "test_data_0600.txt";
test_data_files[601] = "test_data_0601.txt";
test_data_files[602] = "test_data_0602.txt";
test_data_files[603] = "test_data_0603.txt";
test_data_files[604] = "test_data_0604.txt";
test_data_files[605] = "test_data_0605.txt";
test_data_files[606] = "test_data_0606.txt";
test_data_files[607] = "test_data_0607.txt";
test_data_files[608] = "test_data_0608.txt";
test_data_files[609] = "test_data_0609.txt";
test_data_files[610] = "test_data_0610.txt";
test_data_files[611] = "test_data_0611.txt";
test_data_files[612] = "test_data_0612.txt";
test_data_files[613] = "test_data_0613.txt";
test_data_files[614] = "test_data_0614.txt";
test_data_files[615] = "test_data_0615.txt";
test_data_files[616] = "test_data_0616.txt";
test_data_files[617] = "test_data_0617.txt";
test_data_files[618] = "test_data_0618.txt";
test_data_files[619] = "test_data_0619.txt";
test_data_files[620] = "test_data_0620.txt";
test_data_files[621] = "test_data_0621.txt";
test_data_files[622] = "test_data_0622.txt";
test_data_files[623] = "test_data_0623.txt";
test_data_files[624] = "test_data_0624.txt";
test_data_files[625] = "test_data_0625.txt";
test_data_files[626] = "test_data_0626.txt";
test_data_files[627] = "test_data_0627.txt";
test_data_files[628] = "test_data_0628.txt";
test_data_files[629] = "test_data_0629.txt";
test_data_files[630] = "test_data_0630.txt";
test_data_files[631] = "test_data_0631.txt";
test_data_files[632] = "test_data_0632.txt";
test_data_files[633] = "test_data_0633.txt";
test_data_files[634] = "test_data_0634.txt";
test_data_files[635] = "test_data_0635.txt";
test_data_files[636] = "test_data_0636.txt";
test_data_files[637] = "test_data_0637.txt";
test_data_files[638] = "test_data_0638.txt";
test_data_files[639] = "test_data_0639.txt";
test_data_files[640] = "test_data_0640.txt";
test_data_files[641] = "test_data_0641.txt";
test_data_files[642] = "test_data_0642.txt";
test_data_files[643] = "test_data_0643.txt";
test_data_files[644] = "test_data_0644.txt";
test_data_files[645] = "test_data_0645.txt";
test_data_files[646] = "test_data_0646.txt";
test_data_files[647] = "test_data_0647.txt";
test_data_files[648] = "test_data_0648.txt";
test_data_files[649] = "test_data_0649.txt";
test_data_files[650] = "test_data_0650.txt";
test_data_files[651] = "test_data_0651.txt";
test_data_files[652] = "test_data_0652.txt";
test_data_files[653] = "test_data_0653.txt";
test_data_files[654] = "test_data_0654.txt";
test_data_files[655] = "test_data_0655.txt";
test_data_files[656] = "test_data_0656.txt";
test_data_files[657] = "test_data_0657.txt";
test_data_files[658] = "test_data_0658.txt";
test_data_files[659] = "test_data_0659.txt";
test_data_files[660] = "test_data_0660.txt";
test_data_files[661] = "test_data_0661.txt";
test_data_files[662] = "test_data_0662.txt";
test_data_files[663] = "test_data_0663.txt";
test_data_files[664] = "test_data_0664.txt";
test_data_files[665] = "test_data_0665.txt";
test_data_files[666] = "test_data_0666.txt";
test_data_files[667] = "test_data_0667.txt";
test_data_files[668] = "test_data_0668.txt";
test_data_files[669] = "test_data_0669.txt";
test_data_files[670] = "test_data_0670.txt";
test_data_files[671] = "test_data_0671.txt";
test_data_files[672] = "test_data_0672.txt";
test_data_files[673] = "test_data_0673.txt";
test_data_files[674] = "test_data_0674.txt";
test_data_files[675] = "test_data_0675.txt";
test_data_files[676] = "test_data_0676.txt";
test_data_files[677] = "test_data_0677.txt";
test_data_files[678] = "test_data_0678.txt";
test_data_files[679] = "test_data_0679.txt";
test_data_files[680] = "test_data_0680.txt";
test_data_files[681] = "test_data_0681.txt";
test_data_files[682] = "test_data_0682.txt";
test_data_files[683] = "test_data_0683.txt";
test_data_files[684] = "test_data_0684.txt";
test_data_files[685] = "test_data_0685.txt";
test_data_files[686] = "test_data_0686.txt";
test_data_files[687] = "test_data_0687.txt";
test_data_files[688] = "test_data_0688.txt";
test_data_files[689] = "test_data_0689.txt";
test_data_files[690] = "test_data_0690.txt";
test_data_files[691] = "test_data_0691.txt";
test_data_files[692] = "test_data_0692.txt";
test_data_files[693] = "test_data_0693.txt";
test_data_files[694] = "test_data_0694.txt";
test_data_files[695] = "test_data_0695.txt";
test_data_files[696] = "test_data_0696.txt";
test_data_files[697] = "test_data_0697.txt";
test_data_files[698] = "test_data_0698.txt";
test_data_files[699] = "test_data_0699.txt";
test_data_files[700] = "test_data_0700.txt";
test_data_files[701] = "test_data_0701.txt";
test_data_files[702] = "test_data_0702.txt";
test_data_files[703] = "test_data_0703.txt";
test_data_files[704] = "test_data_0704.txt";
test_data_files[705] = "test_data_0705.txt";
test_data_files[706] = "test_data_0706.txt";
test_data_files[707] = "test_data_0707.txt";
test_data_files[708] = "test_data_0708.txt";
test_data_files[709] = "test_data_0709.txt";
test_data_files[710] = "test_data_0710.txt";
test_data_files[711] = "test_data_0711.txt";
test_data_files[712] = "test_data_0712.txt";
test_data_files[713] = "test_data_0713.txt";
test_data_files[714] = "test_data_0714.txt";
test_data_files[715] = "test_data_0715.txt";
test_data_files[716] = "test_data_0716.txt";
test_data_files[717] = "test_data_0717.txt";
test_data_files[718] = "test_data_0718.txt";
test_data_files[719] = "test_data_0719.txt";
test_data_files[720] = "test_data_0720.txt";
test_data_files[721] = "test_data_0721.txt";
test_data_files[722] = "test_data_0722.txt";
test_data_files[723] = "test_data_0723.txt";
test_data_files[724] = "test_data_0724.txt";
test_data_files[725] = "test_data_0725.txt";
test_data_files[726] = "test_data_0726.txt";
test_data_files[727] = "test_data_0727.txt";
test_data_files[728] = "test_data_0728.txt";
test_data_files[729] = "test_data_0729.txt";
test_data_files[730] = "test_data_0730.txt";
test_data_files[731] = "test_data_0731.txt";
test_data_files[732] = "test_data_0732.txt";
test_data_files[733] = "test_data_0733.txt";
test_data_files[734] = "test_data_0734.txt";
test_data_files[735] = "test_data_0735.txt";
test_data_files[736] = "test_data_0736.txt";
test_data_files[737] = "test_data_0737.txt";
test_data_files[738] = "test_data_0738.txt";
test_data_files[739] = "test_data_0739.txt";
test_data_files[740] = "test_data_0740.txt";
test_data_files[741] = "test_data_0741.txt";
test_data_files[742] = "test_data_0742.txt";
test_data_files[743] = "test_data_0743.txt";
test_data_files[744] = "test_data_0744.txt";
test_data_files[745] = "test_data_0745.txt";
test_data_files[746] = "test_data_0746.txt";
test_data_files[747] = "test_data_0747.txt";
test_data_files[748] = "test_data_0748.txt";
test_data_files[749] = "test_data_0749.txt";
test_data_files[750] = "test_data_0750.txt";
test_data_files[751] = "test_data_0751.txt";
test_data_files[752] = "test_data_0752.txt";
test_data_files[753] = "test_data_0753.txt";
test_data_files[754] = "test_data_0754.txt";
test_data_files[755] = "test_data_0755.txt";
test_data_files[756] = "test_data_0756.txt";
test_data_files[757] = "test_data_0757.txt";
test_data_files[758] = "test_data_0758.txt";
test_data_files[759] = "test_data_0759.txt";
test_data_files[760] = "test_data_0760.txt";
test_data_files[761] = "test_data_0761.txt";
test_data_files[762] = "test_data_0762.txt";
test_data_files[763] = "test_data_0763.txt";
test_data_files[764] = "test_data_0764.txt";
test_data_files[765] = "test_data_0765.txt";
test_data_files[766] = "test_data_0766.txt";
test_data_files[767] = "test_data_0767.txt";
test_data_files[768] = "test_data_0768.txt";
test_data_files[769] = "test_data_0769.txt";
test_data_files[770] = "test_data_0770.txt";
test_data_files[771] = "test_data_0771.txt";
test_data_files[772] = "test_data_0772.txt";
test_data_files[773] = "test_data_0773.txt";
test_data_files[774] = "test_data_0774.txt";
test_data_files[775] = "test_data_0775.txt";
test_data_files[776] = "test_data_0776.txt";
test_data_files[777] = "test_data_0777.txt";
test_data_files[778] = "test_data_0778.txt";
test_data_files[779] = "test_data_0779.txt";
test_data_files[780] = "test_data_0780.txt";
test_data_files[781] = "test_data_0781.txt";
test_data_files[782] = "test_data_0782.txt";
test_data_files[783] = "test_data_0783.txt";
test_data_files[784] = "test_data_0784.txt";
test_data_files[785] = "test_data_0785.txt";
test_data_files[786] = "test_data_0786.txt";
test_data_files[787] = "test_data_0787.txt";
test_data_files[788] = "test_data_0788.txt";
test_data_files[789] = "test_data_0789.txt";
test_data_files[790] = "test_data_0790.txt";
test_data_files[791] = "test_data_0791.txt";
test_data_files[792] = "test_data_0792.txt";
test_data_files[793] = "test_data_0793.txt";
test_data_files[794] = "test_data_0794.txt";
test_data_files[795] = "test_data_0795.txt";
test_data_files[796] = "test_data_0796.txt";
test_data_files[797] = "test_data_0797.txt";
test_data_files[798] = "test_data_0798.txt";
test_data_files[799] = "test_data_0799.txt";
test_data_files[800] = "test_data_0800.txt";
test_data_files[801] = "test_data_0801.txt";
test_data_files[802] = "test_data_0802.txt";
test_data_files[803] = "test_data_0803.txt";
test_data_files[804] = "test_data_0804.txt";
test_data_files[805] = "test_data_0805.txt";
test_data_files[806] = "test_data_0806.txt";
test_data_files[807] = "test_data_0807.txt";
test_data_files[808] = "test_data_0808.txt";
test_data_files[809] = "test_data_0809.txt";
test_data_files[810] = "test_data_0810.txt";
test_data_files[811] = "test_data_0811.txt";
test_data_files[812] = "test_data_0812.txt";
test_data_files[813] = "test_data_0813.txt";
test_data_files[814] = "test_data_0814.txt";
test_data_files[815] = "test_data_0815.txt";
test_data_files[816] = "test_data_0816.txt";
test_data_files[817] = "test_data_0817.txt";
test_data_files[818] = "test_data_0818.txt";
test_data_files[819] = "test_data_0819.txt";
test_data_files[820] = "test_data_0820.txt";
test_data_files[821] = "test_data_0821.txt";
test_data_files[822] = "test_data_0822.txt";
test_data_files[823] = "test_data_0823.txt";
test_data_files[824] = "test_data_0824.txt";
test_data_files[825] = "test_data_0825.txt";
test_data_files[826] = "test_data_0826.txt";
test_data_files[827] = "test_data_0827.txt";
test_data_files[828] = "test_data_0828.txt";
test_data_files[829] = "test_data_0829.txt";
test_data_files[830] = "test_data_0830.txt";
test_data_files[831] = "test_data_0831.txt";
test_data_files[832] = "test_data_0832.txt";
test_data_files[833] = "test_data_0833.txt";
test_data_files[834] = "test_data_0834.txt";
test_data_files[835] = "test_data_0835.txt";
test_data_files[836] = "test_data_0836.txt";
test_data_files[837] = "test_data_0837.txt";
test_data_files[838] = "test_data_0838.txt";
test_data_files[839] = "test_data_0839.txt";
test_data_files[840] = "test_data_0840.txt";
test_data_files[841] = "test_data_0841.txt";
test_data_files[842] = "test_data_0842.txt";
test_data_files[843] = "test_data_0843.txt";
test_data_files[844] = "test_data_0844.txt";
test_data_files[845] = "test_data_0845.txt";
test_data_files[846] = "test_data_0846.txt";
test_data_files[847] = "test_data_0847.txt";
test_data_files[848] = "test_data_0848.txt";
test_data_files[849] = "test_data_0849.txt";
test_data_files[850] = "test_data_0850.txt";
test_data_files[851] = "test_data_0851.txt";
test_data_files[852] = "test_data_0852.txt";
test_data_files[853] = "test_data_0853.txt";
test_data_files[854] = "test_data_0854.txt";
test_data_files[855] = "test_data_0855.txt";
test_data_files[856] = "test_data_0856.txt";
test_data_files[857] = "test_data_0857.txt";
test_data_files[858] = "test_data_0858.txt";
test_data_files[859] = "test_data_0859.txt";
test_data_files[860] = "test_data_0860.txt";
test_data_files[861] = "test_data_0861.txt";
test_data_files[862] = "test_data_0862.txt";
test_data_files[863] = "test_data_0863.txt";
test_data_files[864] = "test_data_0864.txt";
test_data_files[865] = "test_data_0865.txt";
test_data_files[866] = "test_data_0866.txt";
test_data_files[867] = "test_data_0867.txt";
test_data_files[868] = "test_data_0868.txt";
test_data_files[869] = "test_data_0869.txt";
test_data_files[870] = "test_data_0870.txt";
test_data_files[871] = "test_data_0871.txt";
test_data_files[872] = "test_data_0872.txt";
test_data_files[873] = "test_data_0873.txt";
test_data_files[874] = "test_data_0874.txt";
test_data_files[875] = "test_data_0875.txt";
test_data_files[876] = "test_data_0876.txt";
test_data_files[877] = "test_data_0877.txt";
test_data_files[878] = "test_data_0878.txt";
test_data_files[879] = "test_data_0879.txt";
test_data_files[880] = "test_data_0880.txt";
test_data_files[881] = "test_data_0881.txt";
test_data_files[882] = "test_data_0882.txt";
test_data_files[883] = "test_data_0883.txt";
test_data_files[884] = "test_data_0884.txt";
test_data_files[885] = "test_data_0885.txt";
test_data_files[886] = "test_data_0886.txt";
test_data_files[887] = "test_data_0887.txt";
test_data_files[888] = "test_data_0888.txt";
test_data_files[889] = "test_data_0889.txt";
test_data_files[890] = "test_data_0890.txt";
test_data_files[891] = "test_data_0891.txt";
test_data_files[892] = "test_data_0892.txt";
test_data_files[893] = "test_data_0893.txt";
test_data_files[894] = "test_data_0894.txt";
test_data_files[895] = "test_data_0895.txt";
test_data_files[896] = "test_data_0896.txt";
test_data_files[897] = "test_data_0897.txt";
test_data_files[898] = "test_data_0898.txt";
test_data_files[899] = "test_data_0899.txt";
test_data_files[900] = "test_data_0900.txt";
test_data_files[901] = "test_data_0901.txt";
test_data_files[902] = "test_data_0902.txt";
test_data_files[903] = "test_data_0903.txt";
test_data_files[904] = "test_data_0904.txt";
test_data_files[905] = "test_data_0905.txt";
test_data_files[906] = "test_data_0906.txt";
test_data_files[907] = "test_data_0907.txt";
test_data_files[908] = "test_data_0908.txt";
test_data_files[909] = "test_data_0909.txt";
test_data_files[910] = "test_data_0910.txt";
test_data_files[911] = "test_data_0911.txt";
test_data_files[912] = "test_data_0912.txt";
test_data_files[913] = "test_data_0913.txt";
test_data_files[914] = "test_data_0914.txt";
test_data_files[915] = "test_data_0915.txt";
test_data_files[916] = "test_data_0916.txt";
test_data_files[917] = "test_data_0917.txt";
test_data_files[918] = "test_data_0918.txt";
test_data_files[919] = "test_data_0919.txt";
test_data_files[920] = "test_data_0920.txt";
test_data_files[921] = "test_data_0921.txt";
test_data_files[922] = "test_data_0922.txt";
test_data_files[923] = "test_data_0923.txt";
test_data_files[924] = "test_data_0924.txt";
test_data_files[925] = "test_data_0925.txt";
test_data_files[926] = "test_data_0926.txt";
test_data_files[927] = "test_data_0927.txt";
test_data_files[928] = "test_data_0928.txt";
test_data_files[929] = "test_data_0929.txt";
test_data_files[930] = "test_data_0930.txt";
test_data_files[931] = "test_data_0931.txt";
test_data_files[932] = "test_data_0932.txt";
test_data_files[933] = "test_data_0933.txt";
test_data_files[934] = "test_data_0934.txt";
test_data_files[935] = "test_data_0935.txt";
test_data_files[936] = "test_data_0936.txt";
test_data_files[937] = "test_data_0937.txt";
test_data_files[938] = "test_data_0938.txt";
test_data_files[939] = "test_data_0939.txt";
test_data_files[940] = "test_data_0940.txt";
test_data_files[941] = "test_data_0941.txt";
test_data_files[942] = "test_data_0942.txt";
test_data_files[943] = "test_data_0943.txt";
test_data_files[944] = "test_data_0944.txt";
test_data_files[945] = "test_data_0945.txt";
test_data_files[946] = "test_data_0946.txt";
test_data_files[947] = "test_data_0947.txt";
test_data_files[948] = "test_data_0948.txt";
test_data_files[949] = "test_data_0949.txt";
test_data_files[950] = "test_data_0950.txt";
test_data_files[951] = "test_data_0951.txt";
test_data_files[952] = "test_data_0952.txt";
test_data_files[953] = "test_data_0953.txt";
test_data_files[954] = "test_data_0954.txt";
test_data_files[955] = "test_data_0955.txt";
test_data_files[956] = "test_data_0956.txt";
test_data_files[957] = "test_data_0957.txt";
test_data_files[958] = "test_data_0958.txt";
test_data_files[959] = "test_data_0959.txt";
test_data_files[960] = "test_data_0960.txt";
test_data_files[961] = "test_data_0961.txt";
test_data_files[962] = "test_data_0962.txt";
test_data_files[963] = "test_data_0963.txt";
test_data_files[964] = "test_data_0964.txt";
test_data_files[965] = "test_data_0965.txt";
test_data_files[966] = "test_data_0966.txt";
test_data_files[967] = "test_data_0967.txt";
test_data_files[968] = "test_data_0968.txt";
test_data_files[969] = "test_data_0969.txt";
test_data_files[970] = "test_data_0970.txt";
test_data_files[971] = "test_data_0971.txt";
test_data_files[972] = "test_data_0972.txt";
test_data_files[973] = "test_data_0973.txt";
test_data_files[974] = "test_data_0974.txt";
test_data_files[975] = "test_data_0975.txt";
test_data_files[976] = "test_data_0976.txt";
test_data_files[977] = "test_data_0977.txt";
test_data_files[978] = "test_data_0978.txt";
test_data_files[979] = "test_data_0979.txt";
test_data_files[980] = "test_data_0980.txt";
test_data_files[981] = "test_data_0981.txt";
test_data_files[982] = "test_data_0982.txt";
test_data_files[983] = "test_data_0983.txt";
test_data_files[984] = "test_data_0984.txt";
test_data_files[985] = "test_data_0985.txt";
test_data_files[986] = "test_data_0986.txt";
test_data_files[987] = "test_data_0987.txt";
test_data_files[988] = "test_data_0988.txt";
test_data_files[989] = "test_data_0989.txt";
test_data_files[990] = "test_data_0990.txt";
test_data_files[991] = "test_data_0991.txt";
test_data_files[992] = "test_data_0992.txt";
test_data_files[993] = "test_data_0993.txt";
test_data_files[994] = "test_data_0994.txt";
test_data_files[995] = "test_data_0995.txt";
test_data_files[996] = "test_data_0996.txt";
test_data_files[997] = "test_data_0997.txt";
test_data_files[998] = "test_data_0998.txt";
test_data_files[999] = "test_data_0999.txt";
test_data_files[1000] = "test_data_1000.txt";
test_data_files[1001] = "test_data_1001.txt";
test_data_files[1002] = "test_data_1002.txt";
test_data_files[1003] = "test_data_1003.txt";
test_data_files[1004] = "test_data_1004.txt";
test_data_files[1005] = "test_data_1005.txt";
test_data_files[1006] = "test_data_1006.txt";
test_data_files[1007] = "test_data_1007.txt";
test_data_files[1008] = "test_data_1008.txt";
test_data_files[1009] = "test_data_1009.txt";
test_data_files[1010] = "test_data_1010.txt";
test_data_files[1011] = "test_data_1011.txt";
test_data_files[1012] = "test_data_1012.txt";
test_data_files[1013] = "test_data_1013.txt";
test_data_files[1014] = "test_data_1014.txt";
test_data_files[1015] = "test_data_1015.txt";
test_data_files[1016] = "test_data_1016.txt";
test_data_files[1017] = "test_data_1017.txt";
test_data_files[1018] = "test_data_1018.txt";
test_data_files[1019] = "test_data_1019.txt";
test_data_files[1020] = "test_data_1020.txt";
test_data_files[1021] = "test_data_1021.txt";
test_data_files[1022] = "test_data_1022.txt";
test_data_files[1023] = "test_data_1023.txt";
test_data_files[1024] = "test_data_1024.txt";
test_data_files[1025] = "test_data_1025.txt";
test_data_files[1026] = "test_data_1026.txt";
test_data_files[1027] = "test_data_1027.txt";
test_data_files[1028] = "test_data_1028.txt";
test_data_files[1029] = "test_data_1029.txt";
test_data_files[1030] = "test_data_1030.txt";
test_data_files[1031] = "test_data_1031.txt";
test_data_files[1032] = "test_data_1032.txt";
test_data_files[1033] = "test_data_1033.txt";
test_data_files[1034] = "test_data_1034.txt";
test_data_files[1035] = "test_data_1035.txt";
test_data_files[1036] = "test_data_1036.txt";
test_data_files[1037] = "test_data_1037.txt";
test_data_files[1038] = "test_data_1038.txt";
test_data_files[1039] = "test_data_1039.txt";
test_data_files[1040] = "test_data_1040.txt";
test_data_files[1041] = "test_data_1041.txt";
test_data_files[1042] = "test_data_1042.txt";
test_data_files[1043] = "test_data_1043.txt";
test_data_files[1044] = "test_data_1044.txt";
test_data_files[1045] = "test_data_1045.txt";
test_data_files[1046] = "test_data_1046.txt";
test_data_files[1047] = "test_data_1047.txt";
test_data_files[1048] = "test_data_1048.txt";
test_data_files[1049] = "test_data_1049.txt";
test_data_files[1050] = "test_data_1050.txt";
test_data_files[1051] = "test_data_1051.txt";
test_data_files[1052] = "test_data_1052.txt";
test_data_files[1053] = "test_data_1053.txt";
test_data_files[1054] = "test_data_1054.txt";
test_data_files[1055] = "test_data_1055.txt";
test_data_files[1056] = "test_data_1056.txt";
test_data_files[1057] = "test_data_1057.txt";
test_data_files[1058] = "test_data_1058.txt";
test_data_files[1059] = "test_data_1059.txt";
test_data_files[1060] = "test_data_1060.txt";
test_data_files[1061] = "test_data_1061.txt";
test_data_files[1062] = "test_data_1062.txt";
test_data_files[1063] = "test_data_1063.txt";
test_data_files[1064] = "test_data_1064.txt";
test_data_files[1065] = "test_data_1065.txt";
test_data_files[1066] = "test_data_1066.txt";
test_data_files[1067] = "test_data_1067.txt";
test_data_files[1068] = "test_data_1068.txt";
test_data_files[1069] = "test_data_1069.txt";
test_data_files[1070] = "test_data_1070.txt";
test_data_files[1071] = "test_data_1071.txt";
test_data_files[1072] = "test_data_1072.txt";
test_data_files[1073] = "test_data_1073.txt";
test_data_files[1074] = "test_data_1074.txt";
test_data_files[1075] = "test_data_1075.txt";
test_data_files[1076] = "test_data_1076.txt";
test_data_files[1077] = "test_data_1077.txt";
test_data_files[1078] = "test_data_1078.txt";
test_data_files[1079] = "test_data_1079.txt";
test_data_files[1080] = "test_data_1080.txt";
test_data_files[1081] = "test_data_1081.txt";
test_data_files[1082] = "test_data_1082.txt";
test_data_files[1083] = "test_data_1083.txt";
test_data_files[1084] = "test_data_1084.txt";
test_data_files[1085] = "test_data_1085.txt";
test_data_files[1086] = "test_data_1086.txt";
test_data_files[1087] = "test_data_1087.txt";
test_data_files[1088] = "test_data_1088.txt";
test_data_files[1089] = "test_data_1089.txt";
test_data_files[1090] = "test_data_1090.txt";
test_data_files[1091] = "test_data_1091.txt";
test_data_files[1092] = "test_data_1092.txt";
test_data_files[1093] = "test_data_1093.txt";
test_data_files[1094] = "test_data_1094.txt";
test_data_files[1095] = "test_data_1095.txt";
test_data_files[1096] = "test_data_1096.txt";
test_data_files[1097] = "test_data_1097.txt";
test_data_files[1098] = "test_data_1098.txt";
test_data_files[1099] = "test_data_1099.txt";
test_data_files[1100] = "test_data_1100.txt";
test_data_files[1101] = "test_data_1101.txt";
test_data_files[1102] = "test_data_1102.txt";
test_data_files[1103] = "test_data_1103.txt";
test_data_files[1104] = "test_data_1104.txt";
test_data_files[1105] = "test_data_1105.txt";
test_data_files[1106] = "test_data_1106.txt";
test_data_files[1107] = "test_data_1107.txt";
test_data_files[1108] = "test_data_1108.txt";
test_data_files[1109] = "test_data_1109.txt";
test_data_files[1110] = "test_data_1110.txt";
test_data_files[1111] = "test_data_1111.txt";
test_data_files[1112] = "test_data_1112.txt";
test_data_files[1113] = "test_data_1113.txt";
test_data_files[1114] = "test_data_1114.txt";
test_data_files[1115] = "test_data_1115.txt";
test_data_files[1116] = "test_data_1116.txt";
test_data_files[1117] = "test_data_1117.txt";
test_data_files[1118] = "test_data_1118.txt";
test_data_files[1119] = "test_data_1119.txt";
test_data_files[1120] = "test_data_1120.txt";
test_data_files[1121] = "test_data_1121.txt";
test_data_files[1122] = "test_data_1122.txt";
test_data_files[1123] = "test_data_1123.txt";
test_data_files[1124] = "test_data_1124.txt";
test_data_files[1125] = "test_data_1125.txt";
test_data_files[1126] = "test_data_1126.txt";
test_data_files[1127] = "test_data_1127.txt";
test_data_files[1128] = "test_data_1128.txt";
test_data_files[1129] = "test_data_1129.txt";
test_data_files[1130] = "test_data_1130.txt";
test_data_files[1131] = "test_data_1131.txt";
test_data_files[1132] = "test_data_1132.txt";
test_data_files[1133] = "test_data_1133.txt";
test_data_files[1134] = "test_data_1134.txt";
test_data_files[1135] = "test_data_1135.txt";
test_data_files[1136] = "test_data_1136.txt";
test_data_files[1137] = "test_data_1137.txt";
test_data_files[1138] = "test_data_1138.txt";
test_data_files[1139] = "test_data_1139.txt";
test_data_files[1140] = "test_data_1140.txt";
test_data_files[1141] = "test_data_1141.txt";
test_data_files[1142] = "test_data_1142.txt";
test_data_files[1143] = "test_data_1143.txt";
test_data_files[1144] = "test_data_1144.txt";
test_data_files[1145] = "test_data_1145.txt";
test_data_files[1146] = "test_data_1146.txt";
test_data_files[1147] = "test_data_1147.txt";
test_data_files[1148] = "test_data_1148.txt";
test_data_files[1149] = "test_data_1149.txt";
test_data_files[1150] = "test_data_1150.txt";
test_data_files[1151] = "test_data_1151.txt";
test_data_files[1152] = "test_data_1152.txt";
test_data_files[1153] = "test_data_1153.txt";
test_data_files[1154] = "test_data_1154.txt";
test_data_files[1155] = "test_data_1155.txt";
test_data_files[1156] = "test_data_1156.txt";
test_data_files[1157] = "test_data_1157.txt";
test_data_files[1158] = "test_data_1158.txt";
test_data_files[1159] = "test_data_1159.txt";
test_data_files[1160] = "test_data_1160.txt";
test_data_files[1161] = "test_data_1161.txt";
test_data_files[1162] = "test_data_1162.txt";
test_data_files[1163] = "test_data_1163.txt";
test_data_files[1164] = "test_data_1164.txt";
test_data_files[1165] = "test_data_1165.txt";
test_data_files[1166] = "test_data_1166.txt";
test_data_files[1167] = "test_data_1167.txt";
test_data_files[1168] = "test_data_1168.txt";
test_data_files[1169] = "test_data_1169.txt";
test_data_files[1170] = "test_data_1170.txt";
test_data_files[1171] = "test_data_1171.txt";
test_data_files[1172] = "test_data_1172.txt";
test_data_files[1173] = "test_data_1173.txt";
test_data_files[1174] = "test_data_1174.txt";
test_data_files[1175] = "test_data_1175.txt";
test_data_files[1176] = "test_data_1176.txt";
test_data_files[1177] = "test_data_1177.txt";
test_data_files[1178] = "test_data_1178.txt";
test_data_files[1179] = "test_data_1179.txt";
test_data_files[1180] = "test_data_1180.txt";
test_data_files[1181] = "test_data_1181.txt";
test_data_files[1182] = "test_data_1182.txt";
test_data_files[1183] = "test_data_1183.txt";
test_data_files[1184] = "test_data_1184.txt";
test_data_files[1185] = "test_data_1185.txt";
test_data_files[1186] = "test_data_1186.txt";
test_data_files[1187] = "test_data_1187.txt";
test_data_files[1188] = "test_data_1188.txt";
test_data_files[1189] = "test_data_1189.txt";
test_data_files[1190] = "test_data_1190.txt";
test_data_files[1191] = "test_data_1191.txt";
test_data_files[1192] = "test_data_1192.txt";
test_data_files[1193] = "test_data_1193.txt";
test_data_files[1194] = "test_data_1194.txt";
test_data_files[1195] = "test_data_1195.txt";
test_data_files[1196] = "test_data_1196.txt";
test_data_files[1197] = "test_data_1197.txt";
test_data_files[1198] = "test_data_1198.txt";
test_data_files[1199] = "test_data_1199.txt";
test_data_files[1200] = "test_data_1200.txt";
test_data_files[1201] = "test_data_1201.txt";
test_data_files[1202] = "test_data_1202.txt";
test_data_files[1203] = "test_data_1203.txt";
test_data_files[1204] = "test_data_1204.txt";
test_data_files[1205] = "test_data_1205.txt";
test_data_files[1206] = "test_data_1206.txt";
test_data_files[1207] = "test_data_1207.txt";
test_data_files[1208] = "test_data_1208.txt";
test_data_files[1209] = "test_data_1209.txt";
test_data_files[1210] = "test_data_1210.txt";
test_data_files[1211] = "test_data_1211.txt";
test_data_files[1212] = "test_data_1212.txt";
test_data_files[1213] = "test_data_1213.txt";
test_data_files[1214] = "test_data_1214.txt";
test_data_files[1215] = "test_data_1215.txt";
test_data_files[1216] = "test_data_1216.txt";
test_data_files[1217] = "test_data_1217.txt";
test_data_files[1218] = "test_data_1218.txt";
test_data_files[1219] = "test_data_1219.txt";
test_data_files[1220] = "test_data_1220.txt";
test_data_files[1221] = "test_data_1221.txt";
test_data_files[1222] = "test_data_1222.txt";
test_data_files[1223] = "test_data_1223.txt";
test_data_files[1224] = "test_data_1224.txt";
test_data_files[1225] = "test_data_1225.txt";
test_data_files[1226] = "test_data_1226.txt";
test_data_files[1227] = "test_data_1227.txt";
test_data_files[1228] = "test_data_1228.txt";
test_data_files[1229] = "test_data_1229.txt";
test_data_files[1230] = "test_data_1230.txt";
test_data_files[1231] = "test_data_1231.txt";
test_data_files[1232] = "test_data_1232.txt";
test_data_files[1233] = "test_data_1233.txt";
test_data_files[1234] = "test_data_1234.txt";
test_data_files[1235] = "test_data_1235.txt";
test_data_files[1236] = "test_data_1236.txt";
test_data_files[1237] = "test_data_1237.txt";
test_data_files[1238] = "test_data_1238.txt";
test_data_files[1239] = "test_data_1239.txt";
test_data_files[1240] = "test_data_1240.txt";
test_data_files[1241] = "test_data_1241.txt";
test_data_files[1242] = "test_data_1242.txt";
test_data_files[1243] = "test_data_1243.txt";
test_data_files[1244] = "test_data_1244.txt";
test_data_files[1245] = "test_data_1245.txt";
test_data_files[1246] = "test_data_1246.txt";
test_data_files[1247] = "test_data_1247.txt";
test_data_files[1248] = "test_data_1248.txt";
test_data_files[1249] = "test_data_1249.txt";
test_data_files[1250] = "test_data_1250.txt";
test_data_files[1251] = "test_data_1251.txt";
test_data_files[1252] = "test_data_1252.txt";
test_data_files[1253] = "test_data_1253.txt";
test_data_files[1254] = "test_data_1254.txt";
test_data_files[1255] = "test_data_1255.txt";
test_data_files[1256] = "test_data_1256.txt";
test_data_files[1257] = "test_data_1257.txt";
test_data_files[1258] = "test_data_1258.txt";
test_data_files[1259] = "test_data_1259.txt";
test_data_files[1260] = "test_data_1260.txt";
test_data_files[1261] = "test_data_1261.txt";
test_data_files[1262] = "test_data_1262.txt";
test_data_files[1263] = "test_data_1263.txt";
test_data_files[1264] = "test_data_1264.txt";
test_data_files[1265] = "test_data_1265.txt";
test_data_files[1266] = "test_data_1266.txt";
test_data_files[1267] = "test_data_1267.txt";
test_data_files[1268] = "test_data_1268.txt";
test_data_files[1269] = "test_data_1269.txt";
test_data_files[1270] = "test_data_1270.txt";
test_data_files[1271] = "test_data_1271.txt";
test_data_files[1272] = "test_data_1272.txt";
test_data_files[1273] = "test_data_1273.txt";
test_data_files[1274] = "test_data_1274.txt";
test_data_files[1275] = "test_data_1275.txt";
test_data_files[1276] = "test_data_1276.txt";
test_data_files[1277] = "test_data_1277.txt";
test_data_files[1278] = "test_data_1278.txt";
test_data_files[1279] = "test_data_1279.txt";
test_data_files[1280] = "test_data_1280.txt";
test_data_files[1281] = "test_data_1281.txt";
test_data_files[1282] = "test_data_1282.txt";
test_data_files[1283] = "test_data_1283.txt";
test_data_files[1284] = "test_data_1284.txt";
test_data_files[1285] = "test_data_1285.txt";
test_data_files[1286] = "test_data_1286.txt";
test_data_files[1287] = "test_data_1287.txt";
test_data_files[1288] = "test_data_1288.txt";
test_data_files[1289] = "test_data_1289.txt";
test_data_files[1290] = "test_data_1290.txt";
test_data_files[1291] = "test_data_1291.txt";
test_data_files[1292] = "test_data_1292.txt";
test_data_files[1293] = "test_data_1293.txt";
test_data_files[1294] = "test_data_1294.txt";
test_data_files[1295] = "test_data_1295.txt";
test_data_files[1296] = "test_data_1296.txt";
test_data_files[1297] = "test_data_1297.txt";
test_data_files[1298] = "test_data_1298.txt";
test_data_files[1299] = "test_data_1299.txt";
test_data_files[1300] = "test_data_1300.txt";
test_data_files[1301] = "test_data_1301.txt";
test_data_files[1302] = "test_data_1302.txt";
test_data_files[1303] = "test_data_1303.txt";
test_data_files[1304] = "test_data_1304.txt";
test_data_files[1305] = "test_data_1305.txt";
test_data_files[1306] = "test_data_1306.txt";
test_data_files[1307] = "test_data_1307.txt";
test_data_files[1308] = "test_data_1308.txt";
test_data_files[1309] = "test_data_1309.txt";
test_data_files[1310] = "test_data_1310.txt";
test_data_files[1311] = "test_data_1311.txt";
test_data_files[1312] = "test_data_1312.txt";
test_data_files[1313] = "test_data_1313.txt";
test_data_files[1314] = "test_data_1314.txt";
test_data_files[1315] = "test_data_1315.txt";
test_data_files[1316] = "test_data_1316.txt";
test_data_files[1317] = "test_data_1317.txt";
test_data_files[1318] = "test_data_1318.txt";
test_data_files[1319] = "test_data_1319.txt";
test_data_files[1320] = "test_data_1320.txt";
test_data_files[1321] = "test_data_1321.txt";
test_data_files[1322] = "test_data_1322.txt";
test_data_files[1323] = "test_data_1323.txt";
test_data_files[1324] = "test_data_1324.txt";
test_data_files[1325] = "test_data_1325.txt";
test_data_files[1326] = "test_data_1326.txt";
test_data_files[1327] = "test_data_1327.txt";
test_data_files[1328] = "test_data_1328.txt";
test_data_files[1329] = "test_data_1329.txt";
test_data_files[1330] = "test_data_1330.txt";
test_data_files[1331] = "test_data_1331.txt";
test_data_files[1332] = "test_data_1332.txt";
test_data_files[1333] = "test_data_1333.txt";
test_data_files[1334] = "test_data_1334.txt";
test_data_files[1335] = "test_data_1335.txt";
test_data_files[1336] = "test_data_1336.txt";
test_data_files[1337] = "test_data_1337.txt";
test_data_files[1338] = "test_data_1338.txt";
test_data_files[1339] = "test_data_1339.txt";
test_data_files[1340] = "test_data_1340.txt";
test_data_files[1341] = "test_data_1341.txt";
test_data_files[1342] = "test_data_1342.txt";
test_data_files[1343] = "test_data_1343.txt";
test_data_files[1344] = "test_data_1344.txt";
test_data_files[1345] = "test_data_1345.txt";
test_data_files[1346] = "test_data_1346.txt";
test_data_files[1347] = "test_data_1347.txt";
test_data_files[1348] = "test_data_1348.txt";
test_data_files[1349] = "test_data_1349.txt";
test_data_files[1350] = "test_data_1350.txt";
test_data_files[1351] = "test_data_1351.txt";
test_data_files[1352] = "test_data_1352.txt";
test_data_files[1353] = "test_data_1353.txt";
test_data_files[1354] = "test_data_1354.txt";
test_data_files[1355] = "test_data_1355.txt";
test_data_files[1356] = "test_data_1356.txt";
test_data_files[1357] = "test_data_1357.txt";
test_data_files[1358] = "test_data_1358.txt";
test_data_files[1359] = "test_data_1359.txt";
test_data_files[1360] = "test_data_1360.txt";
test_data_files[1361] = "test_data_1361.txt";
test_data_files[1362] = "test_data_1362.txt";
test_data_files[1363] = "test_data_1363.txt";
test_data_files[1364] = "test_data_1364.txt";
test_data_files[1365] = "test_data_1365.txt";
test_data_files[1366] = "test_data_1366.txt";
test_data_files[1367] = "test_data_1367.txt";
test_data_files[1368] = "test_data_1368.txt";
test_data_files[1369] = "test_data_1369.txt";
test_data_files[1370] = "test_data_1370.txt";
test_data_files[1371] = "test_data_1371.txt";
test_data_files[1372] = "test_data_1372.txt";
test_data_files[1373] = "test_data_1373.txt";
test_data_files[1374] = "test_data_1374.txt";
test_data_files[1375] = "test_data_1375.txt";
test_data_files[1376] = "test_data_1376.txt";
test_data_files[1377] = "test_data_1377.txt";
test_data_files[1378] = "test_data_1378.txt";
test_data_files[1379] = "test_data_1379.txt";
test_data_files[1380] = "test_data_1380.txt";
test_data_files[1381] = "test_data_1381.txt";
test_data_files[1382] = "test_data_1382.txt";
test_data_files[1383] = "test_data_1383.txt";
test_data_files[1384] = "test_data_1384.txt";
test_data_files[1385] = "test_data_1385.txt";
test_data_files[1386] = "test_data_1386.txt";
test_data_files[1387] = "test_data_1387.txt";
test_data_files[1388] = "test_data_1388.txt";
test_data_files[1389] = "test_data_1389.txt";
test_data_files[1390] = "test_data_1390.txt";
test_data_files[1391] = "test_data_1391.txt";
test_data_files[1392] = "test_data_1392.txt";
test_data_files[1393] = "test_data_1393.txt";
test_data_files[1394] = "test_data_1394.txt";
test_data_files[1395] = "test_data_1395.txt";
test_data_files[1396] = "test_data_1396.txt";
test_data_files[1397] = "test_data_1397.txt";
test_data_files[1398] = "test_data_1398.txt";
test_data_files[1399] = "test_data_1399.txt";
test_data_files[1400] = "test_data_1400.txt";
test_data_files[1401] = "test_data_1401.txt";
test_data_files[1402] = "test_data_1402.txt";
test_data_files[1403] = "test_data_1403.txt";
test_data_files[1404] = "test_data_1404.txt";
test_data_files[1405] = "test_data_1405.txt";
test_data_files[1406] = "test_data_1406.txt";
test_data_files[1407] = "test_data_1407.txt";
test_data_files[1408] = "test_data_1408.txt";
test_data_files[1409] = "test_data_1409.txt";
test_data_files[1410] = "test_data_1410.txt";
test_data_files[1411] = "test_data_1411.txt";
test_data_files[1412] = "test_data_1412.txt";
test_data_files[1413] = "test_data_1413.txt";
test_data_files[1414] = "test_data_1414.txt";
test_data_files[1415] = "test_data_1415.txt";
test_data_files[1416] = "test_data_1416.txt";
test_data_files[1417] = "test_data_1417.txt";
test_data_files[1418] = "test_data_1418.txt";
test_data_files[1419] = "test_data_1419.txt";
test_data_files[1420] = "test_data_1420.txt";
test_data_files[1421] = "test_data_1421.txt";
test_data_files[1422] = "test_data_1422.txt";
test_data_files[1423] = "test_data_1423.txt";
test_data_files[1424] = "test_data_1424.txt";
test_data_files[1425] = "test_data_1425.txt";
test_data_files[1426] = "test_data_1426.txt";
test_data_files[1427] = "test_data_1427.txt";
test_data_files[1428] = "test_data_1428.txt";
test_data_files[1429] = "test_data_1429.txt";
test_data_files[1430] = "test_data_1430.txt";
test_data_files[1431] = "test_data_1431.txt";
test_data_files[1432] = "test_data_1432.txt";
test_data_files[1433] = "test_data_1433.txt";
test_data_files[1434] = "test_data_1434.txt";
test_data_files[1435] = "test_data_1435.txt";
test_data_files[1436] = "test_data_1436.txt";
test_data_files[1437] = "test_data_1437.txt";
test_data_files[1438] = "test_data_1438.txt";
test_data_files[1439] = "test_data_1439.txt";
test_data_files[1440] = "test_data_1440.txt";
test_data_files[1441] = "test_data_1441.txt";
test_data_files[1442] = "test_data_1442.txt";
test_data_files[1443] = "test_data_1443.txt";
test_data_files[1444] = "test_data_1444.txt";
test_data_files[1445] = "test_data_1445.txt";
test_data_files[1446] = "test_data_1446.txt";
test_data_files[1447] = "test_data_1447.txt";
test_data_files[1448] = "test_data_1448.txt";
test_data_files[1449] = "test_data_1449.txt";
test_data_files[1450] = "test_data_1450.txt";
test_data_files[1451] = "test_data_1451.txt";
test_data_files[1452] = "test_data_1452.txt";
test_data_files[1453] = "test_data_1453.txt";
test_data_files[1454] = "test_data_1454.txt";
test_data_files[1455] = "test_data_1455.txt";
test_data_files[1456] = "test_data_1456.txt";
test_data_files[1457] = "test_data_1457.txt";
test_data_files[1458] = "test_data_1458.txt";
test_data_files[1459] = "test_data_1459.txt";
test_data_files[1460] = "test_data_1460.txt";
test_data_files[1461] = "test_data_1461.txt";
test_data_files[1462] = "test_data_1462.txt";
test_data_files[1463] = "test_data_1463.txt";
test_data_files[1464] = "test_data_1464.txt";
test_data_files[1465] = "test_data_1465.txt";
test_data_files[1466] = "test_data_1466.txt";
test_data_files[1467] = "test_data_1467.txt";
test_data_files[1468] = "test_data_1468.txt";
test_data_files[1469] = "test_data_1469.txt";
test_data_files[1470] = "test_data_1470.txt";
test_data_files[1471] = "test_data_1471.txt";
test_data_files[1472] = "test_data_1472.txt";
test_data_files[1473] = "test_data_1473.txt";
test_data_files[1474] = "test_data_1474.txt";
test_data_files[1475] = "test_data_1475.txt";
test_data_files[1476] = "test_data_1476.txt";
test_data_files[1477] = "test_data_1477.txt";
test_data_files[1478] = "test_data_1478.txt";
test_data_files[1479] = "test_data_1479.txt";
test_data_files[1480] = "test_data_1480.txt";
test_data_files[1481] = "test_data_1481.txt";
test_data_files[1482] = "test_data_1482.txt";
test_data_files[1483] = "test_data_1483.txt";
test_data_files[1484] = "test_data_1484.txt";
test_data_files[1485] = "test_data_1485.txt";
test_data_files[1486] = "test_data_1486.txt";
test_data_files[1487] = "test_data_1487.txt";
test_data_files[1488] = "test_data_1488.txt";
test_data_files[1489] = "test_data_1489.txt";
test_data_files[1490] = "test_data_1490.txt";
test_data_files[1491] = "test_data_1491.txt";
test_data_files[1492] = "test_data_1492.txt";
test_data_files[1493] = "test_data_1493.txt";
test_data_files[1494] = "test_data_1494.txt";
test_data_files[1495] = "test_data_1495.txt";
test_data_files[1496] = "test_data_1496.txt";
test_data_files[1497] = "test_data_1497.txt";
test_data_files[1498] = "test_data_1498.txt";
test_data_files[1499] = "test_data_1499.txt";
test_data_files[1500] = "test_data_1500.txt";
test_data_files[1501] = "test_data_1501.txt";
test_data_files[1502] = "test_data_1502.txt";
test_data_files[1503] = "test_data_1503.txt";
test_data_files[1504] = "test_data_1504.txt";
test_data_files[1505] = "test_data_1505.txt";
test_data_files[1506] = "test_data_1506.txt";
test_data_files[1507] = "test_data_1507.txt";
test_data_files[1508] = "test_data_1508.txt";
test_data_files[1509] = "test_data_1509.txt";
test_data_files[1510] = "test_data_1510.txt";
test_data_files[1511] = "test_data_1511.txt";
test_data_files[1512] = "test_data_1512.txt";
test_data_files[1513] = "test_data_1513.txt";
test_data_files[1514] = "test_data_1514.txt";
test_data_files[1515] = "test_data_1515.txt";
test_data_files[1516] = "test_data_1516.txt";
test_data_files[1517] = "test_data_1517.txt";
test_data_files[1518] = "test_data_1518.txt";
test_data_files[1519] = "test_data_1519.txt";
test_data_files[1520] = "test_data_1520.txt";
test_data_files[1521] = "test_data_1521.txt";
test_data_files[1522] = "test_data_1522.txt";
test_data_files[1523] = "test_data_1523.txt";
test_data_files[1524] = "test_data_1524.txt";
test_data_files[1525] = "test_data_1525.txt";
test_data_files[1526] = "test_data_1526.txt";
test_data_files[1527] = "test_data_1527.txt";
test_data_files[1528] = "test_data_1528.txt";
test_data_files[1529] = "test_data_1529.txt";
test_data_files[1530] = "test_data_1530.txt";
test_data_files[1531] = "test_data_1531.txt";
test_data_files[1532] = "test_data_1532.txt";
test_data_files[1533] = "test_data_1533.txt";
test_data_files[1534] = "test_data_1534.txt";
test_data_files[1535] = "test_data_1535.txt";
test_data_files[1536] = "test_data_1536.txt";
test_data_files[1537] = "test_data_1537.txt";
test_data_files[1538] = "test_data_1538.txt";
test_data_files[1539] = "test_data_1539.txt";
test_data_files[1540] = "test_data_1540.txt";
test_data_files[1541] = "test_data_1541.txt";
test_data_files[1542] = "test_data_1542.txt";
test_data_files[1543] = "test_data_1543.txt";
test_data_files[1544] = "test_data_1544.txt";
test_data_files[1545] = "test_data_1545.txt";
test_data_files[1546] = "test_data_1546.txt";
test_data_files[1547] = "test_data_1547.txt";
test_data_files[1548] = "test_data_1548.txt";
test_data_files[1549] = "test_data_1549.txt";
test_data_files[1550] = "test_data_1550.txt";
test_data_files[1551] = "test_data_1551.txt";
test_data_files[1552] = "test_data_1552.txt";
test_data_files[1553] = "test_data_1553.txt";
test_data_files[1554] = "test_data_1554.txt";
test_data_files[1555] = "test_data_1555.txt";
test_data_files[1556] = "test_data_1556.txt";
test_data_files[1557] = "test_data_1557.txt";
test_data_files[1558] = "test_data_1558.txt";
test_data_files[1559] = "test_data_1559.txt";
test_data_files[1560] = "test_data_1560.txt";
test_data_files[1561] = "test_data_1561.txt";
test_data_files[1562] = "test_data_1562.txt";
test_data_files[1563] = "test_data_1563.txt";
test_data_files[1564] = "test_data_1564.txt";
test_data_files[1565] = "test_data_1565.txt";
test_data_files[1566] = "test_data_1566.txt";
test_data_files[1567] = "test_data_1567.txt";
test_data_files[1568] = "test_data_1568.txt";
test_data_files[1569] = "test_data_1569.txt";
test_data_files[1570] = "test_data_1570.txt";
test_data_files[1571] = "test_data_1571.txt";
test_data_files[1572] = "test_data_1572.txt";
test_data_files[1573] = "test_data_1573.txt";
test_data_files[1574] = "test_data_1574.txt";
test_data_files[1575] = "test_data_1575.txt";
test_data_files[1576] = "test_data_1576.txt";
test_data_files[1577] = "test_data_1577.txt";
test_data_files[1578] = "test_data_1578.txt";
test_data_files[1579] = "test_data_1579.txt";
test_data_files[1580] = "test_data_1580.txt";
test_data_files[1581] = "test_data_1581.txt";
test_data_files[1582] = "test_data_1582.txt";
test_data_files[1583] = "test_data_1583.txt";
test_data_files[1584] = "test_data_1584.txt";
test_data_files[1585] = "test_data_1585.txt";
test_data_files[1586] = "test_data_1586.txt";
test_data_files[1587] = "test_data_1587.txt";
test_data_files[1588] = "test_data_1588.txt";
test_data_files[1589] = "test_data_1589.txt";
test_data_files[1590] = "test_data_1590.txt";
test_data_files[1591] = "test_data_1591.txt";
test_data_files[1592] = "test_data_1592.txt";
test_data_files[1593] = "test_data_1593.txt";
test_data_files[1594] = "test_data_1594.txt";
test_data_files[1595] = "test_data_1595.txt";
test_data_files[1596] = "test_data_1596.txt";
test_data_files[1597] = "test_data_1597.txt";
test_data_files[1598] = "test_data_1598.txt";
test_data_files[1599] = "test_data_1599.txt";
test_data_files[1600] = "test_data_1600.txt";
test_data_files[1601] = "test_data_1601.txt";
test_data_files[1602] = "test_data_1602.txt";
test_data_files[1603] = "test_data_1603.txt";
test_data_files[1604] = "test_data_1604.txt";
test_data_files[1605] = "test_data_1605.txt";
test_data_files[1606] = "test_data_1606.txt";
test_data_files[1607] = "test_data_1607.txt";
test_data_files[1608] = "test_data_1608.txt";
test_data_files[1609] = "test_data_1609.txt";
test_data_files[1610] = "test_data_1610.txt";
test_data_files[1611] = "test_data_1611.txt";
test_data_files[1612] = "test_data_1612.txt";
test_data_files[1613] = "test_data_1613.txt";
test_data_files[1614] = "test_data_1614.txt";
test_data_files[1615] = "test_data_1615.txt";
test_data_files[1616] = "test_data_1616.txt";
test_data_files[1617] = "test_data_1617.txt";
test_data_files[1618] = "test_data_1618.txt";
test_data_files[1619] = "test_data_1619.txt";
test_data_files[1620] = "test_data_1620.txt";
test_data_files[1621] = "test_data_1621.txt";
test_data_files[1622] = "test_data_1622.txt";
test_data_files[1623] = "test_data_1623.txt";
test_data_files[1624] = "test_data_1624.txt";
test_data_files[1625] = "test_data_1625.txt";
test_data_files[1626] = "test_data_1626.txt";
test_data_files[1627] = "test_data_1627.txt";
test_data_files[1628] = "test_data_1628.txt";
test_data_files[1629] = "test_data_1629.txt";
test_data_files[1630] = "test_data_1630.txt";
test_data_files[1631] = "test_data_1631.txt";
test_data_files[1632] = "test_data_1632.txt";
test_data_files[1633] = "test_data_1633.txt";
test_data_files[1634] = "test_data_1634.txt";
test_data_files[1635] = "test_data_1635.txt";
test_data_files[1636] = "test_data_1636.txt";
test_data_files[1637] = "test_data_1637.txt";
test_data_files[1638] = "test_data_1638.txt";
test_data_files[1639] = "test_data_1639.txt";
test_data_files[1640] = "test_data_1640.txt";
test_data_files[1641] = "test_data_1641.txt";
test_data_files[1642] = "test_data_1642.txt";
test_data_files[1643] = "test_data_1643.txt";
test_data_files[1644] = "test_data_1644.txt";
test_data_files[1645] = "test_data_1645.txt";
test_data_files[1646] = "test_data_1646.txt";
test_data_files[1647] = "test_data_1647.txt";
test_data_files[1648] = "test_data_1648.txt";
test_data_files[1649] = "test_data_1649.txt";
test_data_files[1650] = "test_data_1650.txt";
test_data_files[1651] = "test_data_1651.txt";
test_data_files[1652] = "test_data_1652.txt";
test_data_files[1653] = "test_data_1653.txt";
test_data_files[1654] = "test_data_1654.txt";
test_data_files[1655] = "test_data_1655.txt";
test_data_files[1656] = "test_data_1656.txt";
test_data_files[1657] = "test_data_1657.txt";
test_data_files[1658] = "test_data_1658.txt";
test_data_files[1659] = "test_data_1659.txt";
test_data_files[1660] = "test_data_1660.txt";
test_data_files[1661] = "test_data_1661.txt";
test_data_files[1662] = "test_data_1662.txt";
test_data_files[1663] = "test_data_1663.txt";
test_data_files[1664] = "test_data_1664.txt";
test_data_files[1665] = "test_data_1665.txt";
test_data_files[1666] = "test_data_1666.txt";
test_data_files[1667] = "test_data_1667.txt";
test_data_files[1668] = "test_data_1668.txt";
test_data_files[1669] = "test_data_1669.txt";
test_data_files[1670] = "test_data_1670.txt";
test_data_files[1671] = "test_data_1671.txt";
test_data_files[1672] = "test_data_1672.txt";
test_data_files[1673] = "test_data_1673.txt";
test_data_files[1674] = "test_data_1674.txt";
test_data_files[1675] = "test_data_1675.txt";
test_data_files[1676] = "test_data_1676.txt";
test_data_files[1677] = "test_data_1677.txt";
test_data_files[1678] = "test_data_1678.txt";
test_data_files[1679] = "test_data_1679.txt";
test_data_files[1680] = "test_data_1680.txt";
test_data_files[1681] = "test_data_1681.txt";
test_data_files[1682] = "test_data_1682.txt";
test_data_files[1683] = "test_data_1683.txt";
test_data_files[1684] = "test_data_1684.txt";
test_data_files[1685] = "test_data_1685.txt";
test_data_files[1686] = "test_data_1686.txt";
test_data_files[1687] = "test_data_1687.txt";
test_data_files[1688] = "test_data_1688.txt";
test_data_files[1689] = "test_data_1689.txt";
test_data_files[1690] = "test_data_1690.txt";
test_data_files[1691] = "test_data_1691.txt";
test_data_files[1692] = "test_data_1692.txt";
test_data_files[1693] = "test_data_1693.txt";
test_data_files[1694] = "test_data_1694.txt";
test_data_files[1695] = "test_data_1695.txt";
test_data_files[1696] = "test_data_1696.txt";
test_data_files[1697] = "test_data_1697.txt";
test_data_files[1698] = "test_data_1698.txt";
test_data_files[1699] = "test_data_1699.txt";
test_data_files[1700] = "test_data_1700.txt";
test_data_files[1701] = "test_data_1701.txt";
test_data_files[1702] = "test_data_1702.txt";
test_data_files[1703] = "test_data_1703.txt";
test_data_files[1704] = "test_data_1704.txt";
test_data_files[1705] = "test_data_1705.txt";
test_data_files[1706] = "test_data_1706.txt";
test_data_files[1707] = "test_data_1707.txt";
test_data_files[1708] = "test_data_1708.txt";
test_data_files[1709] = "test_data_1709.txt";
test_data_files[1710] = "test_data_1710.txt";
test_data_files[1711] = "test_data_1711.txt";
test_data_files[1712] = "test_data_1712.txt";
test_data_files[1713] = "test_data_1713.txt";
test_data_files[1714] = "test_data_1714.txt";
test_data_files[1715] = "test_data_1715.txt";
test_data_files[1716] = "test_data_1716.txt";
test_data_files[1717] = "test_data_1717.txt";
test_data_files[1718] = "test_data_1718.txt";
test_data_files[1719] = "test_data_1719.txt";
test_data_files[1720] = "test_data_1720.txt";
test_data_files[1721] = "test_data_1721.txt";
test_data_files[1722] = "test_data_1722.txt";
test_data_files[1723] = "test_data_1723.txt";
test_data_files[1724] = "test_data_1724.txt";
test_data_files[1725] = "test_data_1725.txt";
test_data_files[1726] = "test_data_1726.txt";
test_data_files[1727] = "test_data_1727.txt";
test_data_files[1728] = "test_data_1728.txt";
test_data_files[1729] = "test_data_1729.txt";
test_data_files[1730] = "test_data_1730.txt";
test_data_files[1731] = "test_data_1731.txt";
test_data_files[1732] = "test_data_1732.txt";
test_data_files[1733] = "test_data_1733.txt";
test_data_files[1734] = "test_data_1734.txt";
test_data_files[1735] = "test_data_1735.txt";
test_data_files[1736] = "test_data_1736.txt";
test_data_files[1737] = "test_data_1737.txt";
test_data_files[1738] = "test_data_1738.txt";
test_data_files[1739] = "test_data_1739.txt";
test_data_files[1740] = "test_data_1740.txt";
test_data_files[1741] = "test_data_1741.txt";
test_data_files[1742] = "test_data_1742.txt";
test_data_files[1743] = "test_data_1743.txt";
test_data_files[1744] = "test_data_1744.txt";
test_data_files[1745] = "test_data_1745.txt";
test_data_files[1746] = "test_data_1746.txt";
test_data_files[1747] = "test_data_1747.txt";
test_data_files[1748] = "test_data_1748.txt";
test_data_files[1749] = "test_data_1749.txt";
test_data_files[1750] = "test_data_1750.txt";
test_data_files[1751] = "test_data_1751.txt";
test_data_files[1752] = "test_data_1752.txt";
test_data_files[1753] = "test_data_1753.txt";
test_data_files[1754] = "test_data_1754.txt";
test_data_files[1755] = "test_data_1755.txt";
test_data_files[1756] = "test_data_1756.txt";
test_data_files[1757] = "test_data_1757.txt";
test_data_files[1758] = "test_data_1758.txt";
test_data_files[1759] = "test_data_1759.txt";
test_data_files[1760] = "test_data_1760.txt";
test_data_files[1761] = "test_data_1761.txt";
test_data_files[1762] = "test_data_1762.txt";
test_data_files[1763] = "test_data_1763.txt";
test_data_files[1764] = "test_data_1764.txt";
test_data_files[1765] = "test_data_1765.txt";
test_data_files[1766] = "test_data_1766.txt";
test_data_files[1767] = "test_data_1767.txt";
test_data_files[1768] = "test_data_1768.txt";
test_data_files[1769] = "test_data_1769.txt";
test_data_files[1770] = "test_data_1770.txt";
test_data_files[1771] = "test_data_1771.txt";
test_data_files[1772] = "test_data_1772.txt";
test_data_files[1773] = "test_data_1773.txt";
test_data_files[1774] = "test_data_1774.txt";
test_data_files[1775] = "test_data_1775.txt";
test_data_files[1776] = "test_data_1776.txt";
test_data_files[1777] = "test_data_1777.txt";
test_data_files[1778] = "test_data_1778.txt";
test_data_files[1779] = "test_data_1779.txt";
test_data_files[1780] = "test_data_1780.txt";
test_data_files[1781] = "test_data_1781.txt";
test_data_files[1782] = "test_data_1782.txt";
test_data_files[1783] = "test_data_1783.txt";
test_data_files[1784] = "test_data_1784.txt";
test_data_files[1785] = "test_data_1785.txt";
test_data_files[1786] = "test_data_1786.txt";
test_data_files[1787] = "test_data_1787.txt";
test_data_files[1788] = "test_data_1788.txt";
test_data_files[1789] = "test_data_1789.txt";
test_data_files[1790] = "test_data_1790.txt";
test_data_files[1791] = "test_data_1791.txt";
test_data_files[1792] = "test_data_1792.txt";
test_data_files[1793] = "test_data_1793.txt";
test_data_files[1794] = "test_data_1794.txt";
test_data_files[1795] = "test_data_1795.txt";
test_data_files[1796] = "test_data_1796.txt";
test_data_files[1797] = "test_data_1797.txt";
test_data_files[1798] = "test_data_1798.txt";
test_data_files[1799] = "test_data_1799.txt";
test_data_files[1800] = "test_data_1800.txt";
test_data_files[1801] = "test_data_1801.txt";
test_data_files[1802] = "test_data_1802.txt";
test_data_files[1803] = "test_data_1803.txt";
test_data_files[1804] = "test_data_1804.txt";
test_data_files[1805] = "test_data_1805.txt";
test_data_files[1806] = "test_data_1806.txt";
test_data_files[1807] = "test_data_1807.txt";
test_data_files[1808] = "test_data_1808.txt";
test_data_files[1809] = "test_data_1809.txt";
test_data_files[1810] = "test_data_1810.txt";
test_data_files[1811] = "test_data_1811.txt";
test_data_files[1812] = "test_data_1812.txt";
test_data_files[1813] = "test_data_1813.txt";
test_data_files[1814] = "test_data_1814.txt";
test_data_files[1815] = "test_data_1815.txt";
test_data_files[1816] = "test_data_1816.txt";
test_data_files[1817] = "test_data_1817.txt";
test_data_files[1818] = "test_data_1818.txt";
test_data_files[1819] = "test_data_1819.txt";
test_data_files[1820] = "test_data_1820.txt";
test_data_files[1821] = "test_data_1821.txt";
test_data_files[1822] = "test_data_1822.txt";
test_data_files[1823] = "test_data_1823.txt";
test_data_files[1824] = "test_data_1824.txt";
test_data_files[1825] = "test_data_1825.txt";
test_data_files[1826] = "test_data_1826.txt";
test_data_files[1827] = "test_data_1827.txt";
test_data_files[1828] = "test_data_1828.txt";
test_data_files[1829] = "test_data_1829.txt";
test_data_files[1830] = "test_data_1830.txt";
test_data_files[1831] = "test_data_1831.txt";
test_data_files[1832] = "test_data_1832.txt";
test_data_files[1833] = "test_data_1833.txt";
test_data_files[1834] = "test_data_1834.txt";
test_data_files[1835] = "test_data_1835.txt";
test_data_files[1836] = "test_data_1836.txt";
test_data_files[1837] = "test_data_1837.txt";
test_data_files[1838] = "test_data_1838.txt";
test_data_files[1839] = "test_data_1839.txt";
test_data_files[1840] = "test_data_1840.txt";
test_data_files[1841] = "test_data_1841.txt";
test_data_files[1842] = "test_data_1842.txt";
test_data_files[1843] = "test_data_1843.txt";
test_data_files[1844] = "test_data_1844.txt";
test_data_files[1845] = "test_data_1845.txt";
test_data_files[1846] = "test_data_1846.txt";
test_data_files[1847] = "test_data_1847.txt";
test_data_files[1848] = "test_data_1848.txt";
test_data_files[1849] = "test_data_1849.txt";
test_data_files[1850] = "test_data_1850.txt";
test_data_files[1851] = "test_data_1851.txt";
test_data_files[1852] = "test_data_1852.txt";
test_data_files[1853] = "test_data_1853.txt";
test_data_files[1854] = "test_data_1854.txt";
test_data_files[1855] = "test_data_1855.txt";
test_data_files[1856] = "test_data_1856.txt";
test_data_files[1857] = "test_data_1857.txt";
test_data_files[1858] = "test_data_1858.txt";
test_data_files[1859] = "test_data_1859.txt";
test_data_files[1860] = "test_data_1860.txt";
test_data_files[1861] = "test_data_1861.txt";
test_data_files[1862] = "test_data_1862.txt";
test_data_files[1863] = "test_data_1863.txt";
test_data_files[1864] = "test_data_1864.txt";
test_data_files[1865] = "test_data_1865.txt";
test_data_files[1866] = "test_data_1866.txt";
test_data_files[1867] = "test_data_1867.txt";
test_data_files[1868] = "test_data_1868.txt";
test_data_files[1869] = "test_data_1869.txt";
test_data_files[1870] = "test_data_1870.txt";
test_data_files[1871] = "test_data_1871.txt";
test_data_files[1872] = "test_data_1872.txt";
test_data_files[1873] = "test_data_1873.txt";
test_data_files[1874] = "test_data_1874.txt";
test_data_files[1875] = "test_data_1875.txt";
test_data_files[1876] = "test_data_1876.txt";
test_data_files[1877] = "test_data_1877.txt";
test_data_files[1878] = "test_data_1878.txt";
test_data_files[1879] = "test_data_1879.txt";
test_data_files[1880] = "test_data_1880.txt";
test_data_files[1881] = "test_data_1881.txt";
test_data_files[1882] = "test_data_1882.txt";
test_data_files[1883] = "test_data_1883.txt";
test_data_files[1884] = "test_data_1884.txt";
test_data_files[1885] = "test_data_1885.txt";
test_data_files[1886] = "test_data_1886.txt";
test_data_files[1887] = "test_data_1887.txt";
test_data_files[1888] = "test_data_1888.txt";
test_data_files[1889] = "test_data_1889.txt";
test_data_files[1890] = "test_data_1890.txt";
test_data_files[1891] = "test_data_1891.txt";
test_data_files[1892] = "test_data_1892.txt";
test_data_files[1893] = "test_data_1893.txt";
test_data_files[1894] = "test_data_1894.txt";
test_data_files[1895] = "test_data_1895.txt";
test_data_files[1896] = "test_data_1896.txt";
test_data_files[1897] = "test_data_1897.txt";
test_data_files[1898] = "test_data_1898.txt";
test_data_files[1899] = "test_data_1899.txt";
test_data_files[1900] = "test_data_1900.txt";
test_data_files[1901] = "test_data_1901.txt";
test_data_files[1902] = "test_data_1902.txt";
test_data_files[1903] = "test_data_1903.txt";
test_data_files[1904] = "test_data_1904.txt";
test_data_files[1905] = "test_data_1905.txt";
test_data_files[1906] = "test_data_1906.txt";
test_data_files[1907] = "test_data_1907.txt";
test_data_files[1908] = "test_data_1908.txt";
test_data_files[1909] = "test_data_1909.txt";
test_data_files[1910] = "test_data_1910.txt";
test_data_files[1911] = "test_data_1911.txt";
test_data_files[1912] = "test_data_1912.txt";
test_data_files[1913] = "test_data_1913.txt";
test_data_files[1914] = "test_data_1914.txt";
test_data_files[1915] = "test_data_1915.txt";
test_data_files[1916] = "test_data_1916.txt";
test_data_files[1917] = "test_data_1917.txt";
test_data_files[1918] = "test_data_1918.txt";
test_data_files[1919] = "test_data_1919.txt";
test_data_files[1920] = "test_data_1920.txt";
test_data_files[1921] = "test_data_1921.txt";
test_data_files[1922] = "test_data_1922.txt";
test_data_files[1923] = "test_data_1923.txt";
test_data_files[1924] = "test_data_1924.txt";
test_data_files[1925] = "test_data_1925.txt";
test_data_files[1926] = "test_data_1926.txt";
test_data_files[1927] = "test_data_1927.txt";
test_data_files[1928] = "test_data_1928.txt";
test_data_files[1929] = "test_data_1929.txt";
test_data_files[1930] = "test_data_1930.txt";
test_data_files[1931] = "test_data_1931.txt";
test_data_files[1932] = "test_data_1932.txt";
test_data_files[1933] = "test_data_1933.txt";
test_data_files[1934] = "test_data_1934.txt";
test_data_files[1935] = "test_data_1935.txt";
test_data_files[1936] = "test_data_1936.txt";
test_data_files[1937] = "test_data_1937.txt";
test_data_files[1938] = "test_data_1938.txt";
test_data_files[1939] = "test_data_1939.txt";
test_data_files[1940] = "test_data_1940.txt";
test_data_files[1941] = "test_data_1941.txt";
test_data_files[1942] = "test_data_1942.txt";
test_data_files[1943] = "test_data_1943.txt";
test_data_files[1944] = "test_data_1944.txt";
test_data_files[1945] = "test_data_1945.txt";
test_data_files[1946] = "test_data_1946.txt";
test_data_files[1947] = "test_data_1947.txt";
test_data_files[1948] = "test_data_1948.txt";
test_data_files[1949] = "test_data_1949.txt";
test_data_files[1950] = "test_data_1950.txt";
test_data_files[1951] = "test_data_1951.txt";
test_data_files[1952] = "test_data_1952.txt";
test_data_files[1953] = "test_data_1953.txt";
test_data_files[1954] = "test_data_1954.txt";
test_data_files[1955] = "test_data_1955.txt";
test_data_files[1956] = "test_data_1956.txt";
test_data_files[1957] = "test_data_1957.txt";
test_data_files[1958] = "test_data_1958.txt";
test_data_files[1959] = "test_data_1959.txt";
test_data_files[1960] = "test_data_1960.txt";
test_data_files[1961] = "test_data_1961.txt";
test_data_files[1962] = "test_data_1962.txt";
test_data_files[1963] = "test_data_1963.txt";
test_data_files[1964] = "test_data_1964.txt";
test_data_files[1965] = "test_data_1965.txt";
test_data_files[1966] = "test_data_1966.txt";
test_data_files[1967] = "test_data_1967.txt";
test_data_files[1968] = "test_data_1968.txt";
test_data_files[1969] = "test_data_1969.txt";
test_data_files[1970] = "test_data_1970.txt";
test_data_files[1971] = "test_data_1971.txt";
test_data_files[1972] = "test_data_1972.txt";
test_data_files[1973] = "test_data_1973.txt";
test_data_files[1974] = "test_data_1974.txt";
test_data_files[1975] = "test_data_1975.txt";
test_data_files[1976] = "test_data_1976.txt";
test_data_files[1977] = "test_data_1977.txt";
test_data_files[1978] = "test_data_1978.txt";
test_data_files[1979] = "test_data_1979.txt";
test_data_files[1980] = "test_data_1980.txt";
test_data_files[1981] = "test_data_1981.txt";
test_data_files[1982] = "test_data_1982.txt";
test_data_files[1983] = "test_data_1983.txt";
test_data_files[1984] = "test_data_1984.txt";
test_data_files[1985] = "test_data_1985.txt";
test_data_files[1986] = "test_data_1986.txt";
test_data_files[1987] = "test_data_1987.txt";
test_data_files[1988] = "test_data_1988.txt";
test_data_files[1989] = "test_data_1989.txt";
test_data_files[1990] = "test_data_1990.txt";
test_data_files[1991] = "test_data_1991.txt";
test_data_files[1992] = "test_data_1992.txt";
test_data_files[1993] = "test_data_1993.txt";
test_data_files[1994] = "test_data_1994.txt";
test_data_files[1995] = "test_data_1995.txt";
test_data_files[1996] = "test_data_1996.txt";
test_data_files[1997] = "test_data_1997.txt";
test_data_files[1998] = "test_data_1998.txt";
test_data_files[1999] = "test_data_1999.txt";
test_data_files[2000] = "test_data_2000.txt";
test_data_files[2001] = "test_data_2001.txt";
test_data_files[2002] = "test_data_2002.txt";
test_data_files[2003] = "test_data_2003.txt";
test_data_files[2004] = "test_data_2004.txt";
test_data_files[2005] = "test_data_2005.txt";
test_data_files[2006] = "test_data_2006.txt";
test_data_files[2007] = "test_data_2007.txt";
test_data_files[2008] = "test_data_2008.txt";
test_data_files[2009] = "test_data_2009.txt";
test_data_files[2010] = "test_data_2010.txt";
test_data_files[2011] = "test_data_2011.txt";
test_data_files[2012] = "test_data_2012.txt";
test_data_files[2013] = "test_data_2013.txt";
test_data_files[2014] = "test_data_2014.txt";
test_data_files[2015] = "test_data_2015.txt";
test_data_files[2016] = "test_data_2016.txt";
test_data_files[2017] = "test_data_2017.txt";
test_data_files[2018] = "test_data_2018.txt";
test_data_files[2019] = "test_data_2019.txt";
test_data_files[2020] = "test_data_2020.txt";
test_data_files[2021] = "test_data_2021.txt";
test_data_files[2022] = "test_data_2022.txt";
test_data_files[2023] = "test_data_2023.txt";
test_data_files[2024] = "test_data_2024.txt";
test_data_files[2025] = "test_data_2025.txt";
test_data_files[2026] = "test_data_2026.txt";
test_data_files[2027] = "test_data_2027.txt";
test_data_files[2028] = "test_data_2028.txt";
test_data_files[2029] = "test_data_2029.txt";
test_data_files[2030] = "test_data_2030.txt";
test_data_files[2031] = "test_data_2031.txt";
test_data_files[2032] = "test_data_2032.txt";
test_data_files[2033] = "test_data_2033.txt";
test_data_files[2034] = "test_data_2034.txt";
test_data_files[2035] = "test_data_2035.txt";
test_data_files[2036] = "test_data_2036.txt";
test_data_files[2037] = "test_data_2037.txt";
test_data_files[2038] = "test_data_2038.txt";
test_data_files[2039] = "test_data_2039.txt";
test_data_files[2040] = "test_data_2040.txt";
test_data_files[2041] = "test_data_2041.txt";
test_data_files[2042] = "test_data_2042.txt";
test_data_files[2043] = "test_data_2043.txt";
test_data_files[2044] = "test_data_2044.txt";
test_data_files[2045] = "test_data_2045.txt";
test_data_files[2046] = "test_data_2046.txt";
test_data_files[2047] = "test_data_2047.txt";
test_data_files[2048] = "test_data_2048.txt";
test_data_files[2049] = "test_data_2049.txt";
test_data_files[2050] = "test_data_2050.txt";
test_data_files[2051] = "test_data_2051.txt";
test_data_files[2052] = "test_data_2052.txt";
test_data_files[2053] = "test_data_2053.txt";
test_data_files[2054] = "test_data_2054.txt";
test_data_files[2055] = "test_data_2055.txt";
test_data_files[2056] = "test_data_2056.txt";
test_data_files[2057] = "test_data_2057.txt";
test_data_files[2058] = "test_data_2058.txt";
test_data_files[2059] = "test_data_2059.txt";
test_data_files[2060] = "test_data_2060.txt";
test_data_files[2061] = "test_data_2061.txt";
test_data_files[2062] = "test_data_2062.txt";
test_data_files[2063] = "test_data_2063.txt";
test_data_files[2064] = "test_data_2064.txt";
test_data_files[2065] = "test_data_2065.txt";
test_data_files[2066] = "test_data_2066.txt";
test_data_files[2067] = "test_data_2067.txt";
test_data_files[2068] = "test_data_2068.txt";
test_data_files[2069] = "test_data_2069.txt";
test_data_files[2070] = "test_data_2070.txt";
test_data_files[2071] = "test_data_2071.txt";
test_data_files[2072] = "test_data_2072.txt";
test_data_files[2073] = "test_data_2073.txt";
test_data_files[2074] = "test_data_2074.txt";
test_data_files[2075] = "test_data_2075.txt";
test_data_files[2076] = "test_data_2076.txt";
test_data_files[2077] = "test_data_2077.txt";
test_data_files[2078] = "test_data_2078.txt";
test_data_files[2079] = "test_data_2079.txt";
test_data_files[2080] = "test_data_2080.txt";
test_data_files[2081] = "test_data_2081.txt";
test_data_files[2082] = "test_data_2082.txt";
test_data_files[2083] = "test_data_2083.txt";
test_data_files[2084] = "test_data_2084.txt";
test_data_files[2085] = "test_data_2085.txt";
test_data_files[2086] = "test_data_2086.txt";
test_data_files[2087] = "test_data_2087.txt";
test_data_files[2088] = "test_data_2088.txt";
test_data_files[2089] = "test_data_2089.txt";
test_data_files[2090] = "test_data_2090.txt";
test_data_files[2091] = "test_data_2091.txt";
test_data_files[2092] = "test_data_2092.txt";
test_data_files[2093] = "test_data_2093.txt";
test_data_files[2094] = "test_data_2094.txt";
test_data_files[2095] = "test_data_2095.txt";
test_data_files[2096] = "test_data_2096.txt";
test_data_files[2097] = "test_data_2097.txt";
test_data_files[2098] = "test_data_2098.txt";
test_data_files[2099] = "test_data_2099.txt";
test_data_files[2100] = "test_data_2100.txt";
test_data_files[2101] = "test_data_2101.txt";
test_data_files[2102] = "test_data_2102.txt";
test_data_files[2103] = "test_data_2103.txt";
test_data_files[2104] = "test_data_2104.txt";
test_data_files[2105] = "test_data_2105.txt";
test_data_files[2106] = "test_data_2106.txt";
test_data_files[2107] = "test_data_2107.txt";
test_data_files[2108] = "test_data_2108.txt";
test_data_files[2109] = "test_data_2109.txt";
test_data_files[2110] = "test_data_2110.txt";
test_data_files[2111] = "test_data_2111.txt";
test_data_files[2112] = "test_data_2112.txt";
test_data_files[2113] = "test_data_2113.txt";
test_data_files[2114] = "test_data_2114.txt";
test_data_files[2115] = "test_data_2115.txt";
test_data_files[2116] = "test_data_2116.txt";
test_data_files[2117] = "test_data_2117.txt";
test_data_files[2118] = "test_data_2118.txt";
test_data_files[2119] = "test_data_2119.txt";
test_data_files[2120] = "test_data_2120.txt";
test_data_files[2121] = "test_data_2121.txt";
test_data_files[2122] = "test_data_2122.txt";
test_data_files[2123] = "test_data_2123.txt";
test_data_files[2124] = "test_data_2124.txt";
test_data_files[2125] = "test_data_2125.txt";
test_data_files[2126] = "test_data_2126.txt";
test_data_files[2127] = "test_data_2127.txt";
test_data_files[2128] = "test_data_2128.txt";
test_data_files[2129] = "test_data_2129.txt";
test_data_files[2130] = "test_data_2130.txt";
test_data_files[2131] = "test_data_2131.txt";
test_data_files[2132] = "test_data_2132.txt";
test_data_files[2133] = "test_data_2133.txt";
test_data_files[2134] = "test_data_2134.txt";
test_data_files[2135] = "test_data_2135.txt";
test_data_files[2136] = "test_data_2136.txt";
test_data_files[2137] = "test_data_2137.txt";
test_data_files[2138] = "test_data_2138.txt";
test_data_files[2139] = "test_data_2139.txt";
test_data_files[2140] = "test_data_2140.txt";
test_data_files[2141] = "test_data_2141.txt";
test_data_files[2142] = "test_data_2142.txt";
test_data_files[2143] = "test_data_2143.txt";
test_data_files[2144] = "test_data_2144.txt";
test_data_files[2145] = "test_data_2145.txt";
test_data_files[2146] = "test_data_2146.txt";
test_data_files[2147] = "test_data_2147.txt";
test_data_files[2148] = "test_data_2148.txt";
test_data_files[2149] = "test_data_2149.txt";
test_data_files[2150] = "test_data_2150.txt";
test_data_files[2151] = "test_data_2151.txt";
test_data_files[2152] = "test_data_2152.txt";
test_data_files[2153] = "test_data_2153.txt";
test_data_files[2154] = "test_data_2154.txt";
test_data_files[2155] = "test_data_2155.txt";
test_data_files[2156] = "test_data_2156.txt";
test_data_files[2157] = "test_data_2157.txt";
test_data_files[2158] = "test_data_2158.txt";
test_data_files[2159] = "test_data_2159.txt";
test_data_files[2160] = "test_data_2160.txt";
test_data_files[2161] = "test_data_2161.txt";
test_data_files[2162] = "test_data_2162.txt";
test_data_files[2163] = "test_data_2163.txt";
test_data_files[2164] = "test_data_2164.txt";
test_data_files[2165] = "test_data_2165.txt";
test_data_files[2166] = "test_data_2166.txt";
test_data_files[2167] = "test_data_2167.txt";
test_data_files[2168] = "test_data_2168.txt";
test_data_files[2169] = "test_data_2169.txt";
test_data_files[2170] = "test_data_2170.txt";
test_data_files[2171] = "test_data_2171.txt";
test_data_files[2172] = "test_data_2172.txt";
test_data_files[2173] = "test_data_2173.txt";
test_data_files[2174] = "test_data_2174.txt";
test_data_files[2175] = "test_data_2175.txt";
test_data_files[2176] = "test_data_2176.txt";
test_data_files[2177] = "test_data_2177.txt";
test_data_files[2178] = "test_data_2178.txt";
test_data_files[2179] = "test_data_2179.txt";
test_data_files[2180] = "test_data_2180.txt";
test_data_files[2181] = "test_data_2181.txt";
test_data_files[2182] = "test_data_2182.txt";
test_data_files[2183] = "test_data_2183.txt";
test_data_files[2184] = "test_data_2184.txt";
test_data_files[2185] = "test_data_2185.txt";
test_data_files[2186] = "test_data_2186.txt";
test_data_files[2187] = "test_data_2187.txt";
test_data_files[2188] = "test_data_2188.txt";
test_data_files[2189] = "test_data_2189.txt";
test_data_files[2190] = "test_data_2190.txt";
test_data_files[2191] = "test_data_2191.txt";
test_data_files[2192] = "test_data_2192.txt";
test_data_files[2193] = "test_data_2193.txt";
test_data_files[2194] = "test_data_2194.txt";
test_data_files[2195] = "test_data_2195.txt";
test_data_files[2196] = "test_data_2196.txt";
test_data_files[2197] = "test_data_2197.txt";
test_data_files[2198] = "test_data_2198.txt";
test_data_files[2199] = "test_data_2199.txt";
test_data_files[2200] = "test_data_2200.txt";
test_data_files[2201] = "test_data_2201.txt";
test_data_files[2202] = "test_data_2202.txt";
test_data_files[2203] = "test_data_2203.txt";
test_data_files[2204] = "test_data_2204.txt";
test_data_files[2205] = "test_data_2205.txt";
test_data_files[2206] = "test_data_2206.txt";
test_data_files[2207] = "test_data_2207.txt";
test_data_files[2208] = "test_data_2208.txt";
test_data_files[2209] = "test_data_2209.txt";
test_data_files[2210] = "test_data_2210.txt";
test_data_files[2211] = "test_data_2211.txt";
test_data_files[2212] = "test_data_2212.txt";
test_data_files[2213] = "test_data_2213.txt";
test_data_files[2214] = "test_data_2214.txt";
test_data_files[2215] = "test_data_2215.txt";
test_data_files[2216] = "test_data_2216.txt";
test_data_files[2217] = "test_data_2217.txt";
test_data_files[2218] = "test_data_2218.txt";
test_data_files[2219] = "test_data_2219.txt";
test_data_files[2220] = "test_data_2220.txt";
test_data_files[2221] = "test_data_2221.txt";
test_data_files[2222] = "test_data_2222.txt";
test_data_files[2223] = "test_data_2223.txt";
test_data_files[2224] = "test_data_2224.txt";
test_data_files[2225] = "test_data_2225.txt";
test_data_files[2226] = "test_data_2226.txt";
test_data_files[2227] = "test_data_2227.txt";
test_data_files[2228] = "test_data_2228.txt";
test_data_files[2229] = "test_data_2229.txt";
test_data_files[2230] = "test_data_2230.txt";
test_data_files[2231] = "test_data_2231.txt";
test_data_files[2232] = "test_data_2232.txt";
test_data_files[2233] = "test_data_2233.txt";
test_data_files[2234] = "test_data_2234.txt";
test_data_files[2235] = "test_data_2235.txt";
test_data_files[2236] = "test_data_2236.txt";
test_data_files[2237] = "test_data_2237.txt";
test_data_files[2238] = "test_data_2238.txt";
test_data_files[2239] = "test_data_2239.txt";
test_data_files[2240] = "test_data_2240.txt";
test_data_files[2241] = "test_data_2241.txt";
test_data_files[2242] = "test_data_2242.txt";
test_data_files[2243] = "test_data_2243.txt";
test_data_files[2244] = "test_data_2244.txt";
test_data_files[2245] = "test_data_2245.txt";
test_data_files[2246] = "test_data_2246.txt";
test_data_files[2247] = "test_data_2247.txt";
test_data_files[2248] = "test_data_2248.txt";
test_data_files[2249] = "test_data_2249.txt";
test_data_files[2250] = "test_data_2250.txt";
test_data_files[2251] = "test_data_2251.txt";
test_data_files[2252] = "test_data_2252.txt";
test_data_files[2253] = "test_data_2253.txt";
test_data_files[2254] = "test_data_2254.txt";
test_data_files[2255] = "test_data_2255.txt";
test_data_files[2256] = "test_data_2256.txt";
test_data_files[2257] = "test_data_2257.txt";
test_data_files[2258] = "test_data_2258.txt";
test_data_files[2259] = "test_data_2259.txt";
test_data_files[2260] = "test_data_2260.txt";
test_data_files[2261] = "test_data_2261.txt";
test_data_files[2262] = "test_data_2262.txt";
test_data_files[2263] = "test_data_2263.txt";
test_data_files[2264] = "test_data_2264.txt";
test_data_files[2265] = "test_data_2265.txt";
test_data_files[2266] = "test_data_2266.txt";
test_data_files[2267] = "test_data_2267.txt";
test_data_files[2268] = "test_data_2268.txt";
test_data_files[2269] = "test_data_2269.txt";
test_data_files[2270] = "test_data_2270.txt";
test_data_files[2271] = "test_data_2271.txt";
test_data_files[2272] = "test_data_2272.txt";
test_data_files[2273] = "test_data_2273.txt";
test_data_files[2274] = "test_data_2274.txt";
test_data_files[2275] = "test_data_2275.txt";
test_data_files[2276] = "test_data_2276.txt";
test_data_files[2277] = "test_data_2277.txt";
test_data_files[2278] = "test_data_2278.txt";
test_data_files[2279] = "test_data_2279.txt";
test_data_files[2280] = "test_data_2280.txt";
test_data_files[2281] = "test_data_2281.txt";
test_data_files[2282] = "test_data_2282.txt";
test_data_files[2283] = "test_data_2283.txt";
test_data_files[2284] = "test_data_2284.txt";
test_data_files[2285] = "test_data_2285.txt";
test_data_files[2286] = "test_data_2286.txt";
test_data_files[2287] = "test_data_2287.txt";
test_data_files[2288] = "test_data_2288.txt";
test_data_files[2289] = "test_data_2289.txt";
test_data_files[2290] = "test_data_2290.txt";
test_data_files[2291] = "test_data_2291.txt";
test_data_files[2292] = "test_data_2292.txt";
test_data_files[2293] = "test_data_2293.txt";
test_data_files[2294] = "test_data_2294.txt";
test_data_files[2295] = "test_data_2295.txt";
test_data_files[2296] = "test_data_2296.txt";
test_data_files[2297] = "test_data_2297.txt";
test_data_files[2298] = "test_data_2298.txt";
test_data_files[2299] = "test_data_2299.txt";
test_data_files[2300] = "test_data_2300.txt";
test_data_files[2301] = "test_data_2301.txt";
test_data_files[2302] = "test_data_2302.txt";
test_data_files[2303] = "test_data_2303.txt";
test_data_files[2304] = "test_data_2304.txt";
test_data_files[2305] = "test_data_2305.txt";
test_data_files[2306] = "test_data_2306.txt";
test_data_files[2307] = "test_data_2307.txt";
test_data_files[2308] = "test_data_2308.txt";
test_data_files[2309] = "test_data_2309.txt";
test_data_files[2310] = "test_data_2310.txt";
test_data_files[2311] = "test_data_2311.txt";
test_data_files[2312] = "test_data_2312.txt";
test_data_files[2313] = "test_data_2313.txt";
test_data_files[2314] = "test_data_2314.txt";
test_data_files[2315] = "test_data_2315.txt";
test_data_files[2316] = "test_data_2316.txt";
test_data_files[2317] = "test_data_2317.txt";
test_data_files[2318] = "test_data_2318.txt";
test_data_files[2319] = "test_data_2319.txt";
test_data_files[2320] = "test_data_2320.txt";
test_data_files[2321] = "test_data_2321.txt";
test_data_files[2322] = "test_data_2322.txt";
test_data_files[2323] = "test_data_2323.txt";
test_data_files[2324] = "test_data_2324.txt";
test_data_files[2325] = "test_data_2325.txt";
test_data_files[2326] = "test_data_2326.txt";
test_data_files[2327] = "test_data_2327.txt";
test_data_files[2328] = "test_data_2328.txt";
test_data_files[2329] = "test_data_2329.txt";
test_data_files[2330] = "test_data_2330.txt";
test_data_files[2331] = "test_data_2331.txt";
test_data_files[2332] = "test_data_2332.txt";
test_data_files[2333] = "test_data_2333.txt";
test_data_files[2334] = "test_data_2334.txt";
test_data_files[2335] = "test_data_2335.txt";
test_data_files[2336] = "test_data_2336.txt";
test_data_files[2337] = "test_data_2337.txt";
test_data_files[2338] = "test_data_2338.txt";
test_data_files[2339] = "test_data_2339.txt";
test_data_files[2340] = "test_data_2340.txt";
test_data_files[2341] = "test_data_2341.txt";
test_data_files[2342] = "test_data_2342.txt";
test_data_files[2343] = "test_data_2343.txt";
test_data_files[2344] = "test_data_2344.txt";
test_data_files[2345] = "test_data_2345.txt";
test_data_files[2346] = "test_data_2346.txt";
test_data_files[2347] = "test_data_2347.txt";
test_data_files[2348] = "test_data_2348.txt";
test_data_files[2349] = "test_data_2349.txt";
test_data_files[2350] = "test_data_2350.txt";
test_data_files[2351] = "test_data_2351.txt";
test_data_files[2352] = "test_data_2352.txt";
test_data_files[2353] = "test_data_2353.txt";
test_data_files[2354] = "test_data_2354.txt";
test_data_files[2355] = "test_data_2355.txt";
test_data_files[2356] = "test_data_2356.txt";
test_data_files[2357] = "test_data_2357.txt";
test_data_files[2358] = "test_data_2358.txt";
test_data_files[2359] = "test_data_2359.txt";
test_data_files[2360] = "test_data_2360.txt";
test_data_files[2361] = "test_data_2361.txt";
test_data_files[2362] = "test_data_2362.txt";
test_data_files[2363] = "test_data_2363.txt";
test_data_files[2364] = "test_data_2364.txt";
test_data_files[2365] = "test_data_2365.txt";
test_data_files[2366] = "test_data_2366.txt";
test_data_files[2367] = "test_data_2367.txt";
test_data_files[2368] = "test_data_2368.txt";
test_data_files[2369] = "test_data_2369.txt";
test_data_files[2370] = "test_data_2370.txt";
test_data_files[2371] = "test_data_2371.txt";
test_data_files[2372] = "test_data_2372.txt";
test_data_files[2373] = "test_data_2373.txt";
test_data_files[2374] = "test_data_2374.txt";
test_data_files[2375] = "test_data_2375.txt";
test_data_files[2376] = "test_data_2376.txt";
test_data_files[2377] = "test_data_2377.txt";
test_data_files[2378] = "test_data_2378.txt";
test_data_files[2379] = "test_data_2379.txt";
test_data_files[2380] = "test_data_2380.txt";
test_data_files[2381] = "test_data_2381.txt";
test_data_files[2382] = "test_data_2382.txt";
test_data_files[2383] = "test_data_2383.txt";
test_data_files[2384] = "test_data_2384.txt";
test_data_files[2385] = "test_data_2385.txt";
test_data_files[2386] = "test_data_2386.txt";
test_data_files[2387] = "test_data_2387.txt";
test_data_files[2388] = "test_data_2388.txt";
test_data_files[2389] = "test_data_2389.txt";
test_data_files[2390] = "test_data_2390.txt";
test_data_files[2391] = "test_data_2391.txt";
test_data_files[2392] = "test_data_2392.txt";
test_data_files[2393] = "test_data_2393.txt";
test_data_files[2394] = "test_data_2394.txt";
test_data_files[2395] = "test_data_2395.txt";
test_data_files[2396] = "test_data_2396.txt";
test_data_files[2397] = "test_data_2397.txt";
test_data_files[2398] = "test_data_2398.txt";
test_data_files[2399] = "test_data_2399.txt";
test_data_files[2400] = "test_data_2400.txt";
test_data_files[2401] = "test_data_2401.txt";
test_data_files[2402] = "test_data_2402.txt";
test_data_files[2403] = "test_data_2403.txt";
test_data_files[2404] = "test_data_2404.txt";
test_data_files[2405] = "test_data_2405.txt";
test_data_files[2406] = "test_data_2406.txt";
test_data_files[2407] = "test_data_2407.txt";
test_data_files[2408] = "test_data_2408.txt";
test_data_files[2409] = "test_data_2409.txt";
test_data_files[2410] = "test_data_2410.txt";
test_data_files[2411] = "test_data_2411.txt";
test_data_files[2412] = "test_data_2412.txt";
test_data_files[2413] = "test_data_2413.txt";
test_data_files[2414] = "test_data_2414.txt";
test_data_files[2415] = "test_data_2415.txt";
test_data_files[2416] = "test_data_2416.txt";
test_data_files[2417] = "test_data_2417.txt";
test_data_files[2418] = "test_data_2418.txt";
test_data_files[2419] = "test_data_2419.txt";
test_data_files[2420] = "test_data_2420.txt";
test_data_files[2421] = "test_data_2421.txt";
test_data_files[2422] = "test_data_2422.txt";
test_data_files[2423] = "test_data_2423.txt";
test_data_files[2424] = "test_data_2424.txt";
test_data_files[2425] = "test_data_2425.txt";
test_data_files[2426] = "test_data_2426.txt";
test_data_files[2427] = "test_data_2427.txt";
test_data_files[2428] = "test_data_2428.txt";
test_data_files[2429] = "test_data_2429.txt";
test_data_files[2430] = "test_data_2430.txt";
test_data_files[2431] = "test_data_2431.txt";
test_data_files[2432] = "test_data_2432.txt";
test_data_files[2433] = "test_data_2433.txt";
test_data_files[2434] = "test_data_2434.txt";
test_data_files[2435] = "test_data_2435.txt";
test_data_files[2436] = "test_data_2436.txt";
test_data_files[2437] = "test_data_2437.txt";
test_data_files[2438] = "test_data_2438.txt";
test_data_files[2439] = "test_data_2439.txt";
test_data_files[2440] = "test_data_2440.txt";
test_data_files[2441] = "test_data_2441.txt";
test_data_files[2442] = "test_data_2442.txt";
test_data_files[2443] = "test_data_2443.txt";
test_data_files[2444] = "test_data_2444.txt";
test_data_files[2445] = "test_data_2445.txt";
test_data_files[2446] = "test_data_2446.txt";
test_data_files[2447] = "test_data_2447.txt";
test_data_files[2448] = "test_data_2448.txt";
test_data_files[2449] = "test_data_2449.txt";
test_data_files[2450] = "test_data_2450.txt";
test_data_files[2451] = "test_data_2451.txt";
test_data_files[2452] = "test_data_2452.txt";
test_data_files[2453] = "test_data_2453.txt";
test_data_files[2454] = "test_data_2454.txt";
test_data_files[2455] = "test_data_2455.txt";
test_data_files[2456] = "test_data_2456.txt";
test_data_files[2457] = "test_data_2457.txt";
test_data_files[2458] = "test_data_2458.txt";
test_data_files[2459] = "test_data_2459.txt";
test_data_files[2460] = "test_data_2460.txt";
test_data_files[2461] = "test_data_2461.txt";
test_data_files[2462] = "test_data_2462.txt";
test_data_files[2463] = "test_data_2463.txt";
test_data_files[2464] = "test_data_2464.txt";
test_data_files[2465] = "test_data_2465.txt";
test_data_files[2466] = "test_data_2466.txt";
test_data_files[2467] = "test_data_2467.txt";
test_data_files[2468] = "test_data_2468.txt";
test_data_files[2469] = "test_data_2469.txt";
test_data_files[2470] = "test_data_2470.txt";
test_data_files[2471] = "test_data_2471.txt";
test_data_files[2472] = "test_data_2472.txt";
test_data_files[2473] = "test_data_2473.txt";
test_data_files[2474] = "test_data_2474.txt";
test_data_files[2475] = "test_data_2475.txt";
test_data_files[2476] = "test_data_2476.txt";
test_data_files[2477] = "test_data_2477.txt";
test_data_files[2478] = "test_data_2478.txt";
test_data_files[2479] = "test_data_2479.txt";
test_data_files[2480] = "test_data_2480.txt";
test_data_files[2481] = "test_data_2481.txt";
test_data_files[2482] = "test_data_2482.txt";
test_data_files[2483] = "test_data_2483.txt";
test_data_files[2484] = "test_data_2484.txt";
test_data_files[2485] = "test_data_2485.txt";
test_data_files[2486] = "test_data_2486.txt";
test_data_files[2487] = "test_data_2487.txt";
test_data_files[2488] = "test_data_2488.txt";
test_data_files[2489] = "test_data_2489.txt";
test_data_files[2490] = "test_data_2490.txt";
test_data_files[2491] = "test_data_2491.txt";
test_data_files[2492] = "test_data_2492.txt";
test_data_files[2493] = "test_data_2493.txt";
test_data_files[2494] = "test_data_2494.txt";
test_data_files[2495] = "test_data_2495.txt";
test_data_files[2496] = "test_data_2496.txt";
test_data_files[2497] = "test_data_2497.txt";
test_data_files[2498] = "test_data_2498.txt";
test_data_files[2499] = "test_data_2499.txt";
test_data_files[2500] = "test_data_2500.txt";
test_data_files[2501] = "test_data_2501.txt";
test_data_files[2502] = "test_data_2502.txt";
test_data_files[2503] = "test_data_2503.txt";
test_data_files[2504] = "test_data_2504.txt";
test_data_files[2505] = "test_data_2505.txt";
test_data_files[2506] = "test_data_2506.txt";
test_data_files[2507] = "test_data_2507.txt";
test_data_files[2508] = "test_data_2508.txt";
test_data_files[2509] = "test_data_2509.txt";
test_data_files[2510] = "test_data_2510.txt";
test_data_files[2511] = "test_data_2511.txt";
test_data_files[2512] = "test_data_2512.txt";
test_data_files[2513] = "test_data_2513.txt";
test_data_files[2514] = "test_data_2514.txt";
test_data_files[2515] = "test_data_2515.txt";
test_data_files[2516] = "test_data_2516.txt";
test_data_files[2517] = "test_data_2517.txt";
test_data_files[2518] = "test_data_2518.txt";
test_data_files[2519] = "test_data_2519.txt";
test_data_files[2520] = "test_data_2520.txt";
test_data_files[2521] = "test_data_2521.txt";
test_data_files[2522] = "test_data_2522.txt";
test_data_files[2523] = "test_data_2523.txt";
test_data_files[2524] = "test_data_2524.txt";
test_data_files[2525] = "test_data_2525.txt";
test_data_files[2526] = "test_data_2526.txt";
test_data_files[2527] = "test_data_2527.txt";
test_data_files[2528] = "test_data_2528.txt";
test_data_files[2529] = "test_data_2529.txt";
test_data_files[2530] = "test_data_2530.txt";
test_data_files[2531] = "test_data_2531.txt";
test_data_files[2532] = "test_data_2532.txt";
test_data_files[2533] = "test_data_2533.txt";
test_data_files[2534] = "test_data_2534.txt";
test_data_files[2535] = "test_data_2535.txt";
test_data_files[2536] = "test_data_2536.txt";
test_data_files[2537] = "test_data_2537.txt";
test_data_files[2538] = "test_data_2538.txt";
test_data_files[2539] = "test_data_2539.txt";
test_data_files[2540] = "test_data_2540.txt";
test_data_files[2541] = "test_data_2541.txt";
test_data_files[2542] = "test_data_2542.txt";
test_data_files[2543] = "test_data_2543.txt";
test_data_files[2544] = "test_data_2544.txt";
test_data_files[2545] = "test_data_2545.txt";
test_data_files[2546] = "test_data_2546.txt";
test_data_files[2547] = "test_data_2547.txt";
test_data_files[2548] = "test_data_2548.txt";
test_data_files[2549] = "test_data_2549.txt";
test_data_files[2550] = "test_data_2550.txt";
test_data_files[2551] = "test_data_2551.txt";
test_data_files[2552] = "test_data_2552.txt";
test_data_files[2553] = "test_data_2553.txt";
test_data_files[2554] = "test_data_2554.txt";
test_data_files[2555] = "test_data_2555.txt";
test_data_files[2556] = "test_data_2556.txt";
test_data_files[2557] = "test_data_2557.txt";
test_data_files[2558] = "test_data_2558.txt";
test_data_files[2559] = "test_data_2559.txt";
test_data_files[2560] = "test_data_2560.txt";
test_data_files[2561] = "test_data_2561.txt";
test_data_files[2562] = "test_data_2562.txt";
test_data_files[2563] = "test_data_2563.txt";
test_data_files[2564] = "test_data_2564.txt";
test_data_files[2565] = "test_data_2565.txt";
test_data_files[2566] = "test_data_2566.txt";
test_data_files[2567] = "test_data_2567.txt";
test_data_files[2568] = "test_data_2568.txt";
test_data_files[2569] = "test_data_2569.txt";
test_data_files[2570] = "test_data_2570.txt";
test_data_files[2571] = "test_data_2571.txt";
test_data_files[2572] = "test_data_2572.txt";
test_data_files[2573] = "test_data_2573.txt";
test_data_files[2574] = "test_data_2574.txt";
test_data_files[2575] = "test_data_2575.txt";
test_data_files[2576] = "test_data_2576.txt";
test_data_files[2577] = "test_data_2577.txt";
test_data_files[2578] = "test_data_2578.txt";
test_data_files[2579] = "test_data_2579.txt";
test_data_files[2580] = "test_data_2580.txt";
test_data_files[2581] = "test_data_2581.txt";
test_data_files[2582] = "test_data_2582.txt";
test_data_files[2583] = "test_data_2583.txt";
test_data_files[2584] = "test_data_2584.txt";
test_data_files[2585] = "test_data_2585.txt";
test_data_files[2586] = "test_data_2586.txt";
test_data_files[2587] = "test_data_2587.txt";
test_data_files[2588] = "test_data_2588.txt";
test_data_files[2589] = "test_data_2589.txt";
test_data_files[2590] = "test_data_2590.txt";
test_data_files[2591] = "test_data_2591.txt";
test_data_files[2592] = "test_data_2592.txt";
test_data_files[2593] = "test_data_2593.txt";
test_data_files[2594] = "test_data_2594.txt";
test_data_files[2595] = "test_data_2595.txt";
test_data_files[2596] = "test_data_2596.txt";
test_data_files[2597] = "test_data_2597.txt";
test_data_files[2598] = "test_data_2598.txt";
test_data_files[2599] = "test_data_2599.txt";
test_data_files[2600] = "test_data_2600.txt";
test_data_files[2601] = "test_data_2601.txt";
test_data_files[2602] = "test_data_2602.txt";
test_data_files[2603] = "test_data_2603.txt";
test_data_files[2604] = "test_data_2604.txt";
test_data_files[2605] = "test_data_2605.txt";
test_data_files[2606] = "test_data_2606.txt";
test_data_files[2607] = "test_data_2607.txt";
test_data_files[2608] = "test_data_2608.txt";
test_data_files[2609] = "test_data_2609.txt";
test_data_files[2610] = "test_data_2610.txt";
test_data_files[2611] = "test_data_2611.txt";
test_data_files[2612] = "test_data_2612.txt";
test_data_files[2613] = "test_data_2613.txt";
test_data_files[2614] = "test_data_2614.txt";
test_data_files[2615] = "test_data_2615.txt";
test_data_files[2616] = "test_data_2616.txt";
test_data_files[2617] = "test_data_2617.txt";
test_data_files[2618] = "test_data_2618.txt";
test_data_files[2619] = "test_data_2619.txt";
test_data_files[2620] = "test_data_2620.txt";
test_data_files[2621] = "test_data_2621.txt";
test_data_files[2622] = "test_data_2622.txt";
test_data_files[2623] = "test_data_2623.txt";
test_data_files[2624] = "test_data_2624.txt";
test_data_files[2625] = "test_data_2625.txt";
test_data_files[2626] = "test_data_2626.txt";
test_data_files[2627] = "test_data_2627.txt";
test_data_files[2628] = "test_data_2628.txt";
test_data_files[2629] = "test_data_2629.txt";
test_data_files[2630] = "test_data_2630.txt";
test_data_files[2631] = "test_data_2631.txt";
test_data_files[2632] = "test_data_2632.txt";
test_data_files[2633] = "test_data_2633.txt";
test_data_files[2634] = "test_data_2634.txt";
test_data_files[2635] = "test_data_2635.txt";
test_data_files[2636] = "test_data_2636.txt";
test_data_files[2637] = "test_data_2637.txt";
test_data_files[2638] = "test_data_2638.txt";
test_data_files[2639] = "test_data_2639.txt";
test_data_files[2640] = "test_data_2640.txt";
test_data_files[2641] = "test_data_2641.txt";
test_data_files[2642] = "test_data_2642.txt";
test_data_files[2643] = "test_data_2643.txt";
test_data_files[2644] = "test_data_2644.txt";
test_data_files[2645] = "test_data_2645.txt";
test_data_files[2646] = "test_data_2646.txt";
test_data_files[2647] = "test_data_2647.txt";
test_data_files[2648] = "test_data_2648.txt";
test_data_files[2649] = "test_data_2649.txt";
test_data_files[2650] = "test_data_2650.txt";
test_data_files[2651] = "test_data_2651.txt";
test_data_files[2652] = "test_data_2652.txt";
test_data_files[2653] = "test_data_2653.txt";
test_data_files[2654] = "test_data_2654.txt";
test_data_files[2655] = "test_data_2655.txt";
test_data_files[2656] = "test_data_2656.txt";
test_data_files[2657] = "test_data_2657.txt";
test_data_files[2658] = "test_data_2658.txt";
test_data_files[2659] = "test_data_2659.txt";
test_data_files[2660] = "test_data_2660.txt";
test_data_files[2661] = "test_data_2661.txt";
test_data_files[2662] = "test_data_2662.txt";
test_data_files[2663] = "test_data_2663.txt";
test_data_files[2664] = "test_data_2664.txt";
test_data_files[2665] = "test_data_2665.txt";
test_data_files[2666] = "test_data_2666.txt";
test_data_files[2667] = "test_data_2667.txt";
test_data_files[2668] = "test_data_2668.txt";
test_data_files[2669] = "test_data_2669.txt";
test_data_files[2670] = "test_data_2670.txt";
test_data_files[2671] = "test_data_2671.txt";
test_data_files[2672] = "test_data_2672.txt";
test_data_files[2673] = "test_data_2673.txt";
test_data_files[2674] = "test_data_2674.txt";
test_data_files[2675] = "test_data_2675.txt";
test_data_files[2676] = "test_data_2676.txt";
test_data_files[2677] = "test_data_2677.txt";
test_data_files[2678] = "test_data_2678.txt";
test_data_files[2679] = "test_data_2679.txt";
test_data_files[2680] = "test_data_2680.txt";
test_data_files[2681] = "test_data_2681.txt";
test_data_files[2682] = "test_data_2682.txt";
test_data_files[2683] = "test_data_2683.txt";
test_data_files[2684] = "test_data_2684.txt";
test_data_files[2685] = "test_data_2685.txt";
test_data_files[2686] = "test_data_2686.txt";
test_data_files[2687] = "test_data_2687.txt";
test_data_files[2688] = "test_data_2688.txt";
test_data_files[2689] = "test_data_2689.txt";
test_data_files[2690] = "test_data_2690.txt";
test_data_files[2691] = "test_data_2691.txt";
test_data_files[2692] = "test_data_2692.txt";
test_data_files[2693] = "test_data_2693.txt";
test_data_files[2694] = "test_data_2694.txt";
test_data_files[2695] = "test_data_2695.txt";
test_data_files[2696] = "test_data_2696.txt";
test_data_files[2697] = "test_data_2697.txt";
test_data_files[2698] = "test_data_2698.txt";
test_data_files[2699] = "test_data_2699.txt";
test_data_files[2700] = "test_data_2700.txt";
test_data_files[2701] = "test_data_2701.txt";
test_data_files[2702] = "test_data_2702.txt";
test_data_files[2703] = "test_data_2703.txt";
test_data_files[2704] = "test_data_2704.txt";
test_data_files[2705] = "test_data_2705.txt";
test_data_files[2706] = "test_data_2706.txt";
test_data_files[2707] = "test_data_2707.txt";
test_data_files[2708] = "test_data_2708.txt";
test_data_files[2709] = "test_data_2709.txt";
test_data_files[2710] = "test_data_2710.txt";
test_data_files[2711] = "test_data_2711.txt";
test_data_files[2712] = "test_data_2712.txt";
test_data_files[2713] = "test_data_2713.txt";
test_data_files[2714] = "test_data_2714.txt";
test_data_files[2715] = "test_data_2715.txt";
test_data_files[2716] = "test_data_2716.txt";
test_data_files[2717] = "test_data_2717.txt";
test_data_files[2718] = "test_data_2718.txt";
test_data_files[2719] = "test_data_2719.txt";
test_data_files[2720] = "test_data_2720.txt";
test_data_files[2721] = "test_data_2721.txt";
test_data_files[2722] = "test_data_2722.txt";
test_data_files[2723] = "test_data_2723.txt";
test_data_files[2724] = "test_data_2724.txt";
test_data_files[2725] = "test_data_2725.txt";
test_data_files[2726] = "test_data_2726.txt";
test_data_files[2727] = "test_data_2727.txt";
test_data_files[2728] = "test_data_2728.txt";
test_data_files[2729] = "test_data_2729.txt";
test_data_files[2730] = "test_data_2730.txt";
test_data_files[2731] = "test_data_2731.txt";
test_data_files[2732] = "test_data_2732.txt";
test_data_files[2733] = "test_data_2733.txt";
test_data_files[2734] = "test_data_2734.txt";
test_data_files[2735] = "test_data_2735.txt";
test_data_files[2736] = "test_data_2736.txt";
test_data_files[2737] = "test_data_2737.txt";
test_data_files[2738] = "test_data_2738.txt";
test_data_files[2739] = "test_data_2739.txt";
test_data_files[2740] = "test_data_2740.txt";
test_data_files[2741] = "test_data_2741.txt";
test_data_files[2742] = "test_data_2742.txt";
test_data_files[2743] = "test_data_2743.txt";
test_data_files[2744] = "test_data_2744.txt";
test_data_files[2745] = "test_data_2745.txt";
test_data_files[2746] = "test_data_2746.txt";
test_data_files[2747] = "test_data_2747.txt";
test_data_files[2748] = "test_data_2748.txt";
test_data_files[2749] = "test_data_2749.txt";
test_data_files[2750] = "test_data_2750.txt";
test_data_files[2751] = "test_data_2751.txt";
test_data_files[2752] = "test_data_2752.txt";
test_data_files[2753] = "test_data_2753.txt";
test_data_files[2754] = "test_data_2754.txt";
test_data_files[2755] = "test_data_2755.txt";
test_data_files[2756] = "test_data_2756.txt";
test_data_files[2757] = "test_data_2757.txt";
test_data_files[2758] = "test_data_2758.txt";
test_data_files[2759] = "test_data_2759.txt";
test_data_files[2760] = "test_data_2760.txt";
test_data_files[2761] = "test_data_2761.txt";
test_data_files[2762] = "test_data_2762.txt";
test_data_files[2763] = "test_data_2763.txt";
test_data_files[2764] = "test_data_2764.txt";
test_data_files[2765] = "test_data_2765.txt";
test_data_files[2766] = "test_data_2766.txt";
test_data_files[2767] = "test_data_2767.txt";
test_data_files[2768] = "test_data_2768.txt";
test_data_files[2769] = "test_data_2769.txt";
test_data_files[2770] = "test_data_2770.txt";
test_data_files[2771] = "test_data_2771.txt";
test_data_files[2772] = "test_data_2772.txt";
test_data_files[2773] = "test_data_2773.txt";
test_data_files[2774] = "test_data_2774.txt";
test_data_files[2775] = "test_data_2775.txt";
test_data_files[2776] = "test_data_2776.txt";
test_data_files[2777] = "test_data_2777.txt";
test_data_files[2778] = "test_data_2778.txt";
test_data_files[2779] = "test_data_2779.txt";
test_data_files[2780] = "test_data_2780.txt";
test_data_files[2781] = "test_data_2781.txt";
test_data_files[2782] = "test_data_2782.txt";
test_data_files[2783] = "test_data_2783.txt";
test_data_files[2784] = "test_data_2784.txt";
test_data_files[2785] = "test_data_2785.txt";
test_data_files[2786] = "test_data_2786.txt";
test_data_files[2787] = "test_data_2787.txt";
test_data_files[2788] = "test_data_2788.txt";
test_data_files[2789] = "test_data_2789.txt";
test_data_files[2790] = "test_data_2790.txt";
test_data_files[2791] = "test_data_2791.txt";
test_data_files[2792] = "test_data_2792.txt";
test_data_files[2793] = "test_data_2793.txt";
test_data_files[2794] = "test_data_2794.txt";
test_data_files[2795] = "test_data_2795.txt";
test_data_files[2796] = "test_data_2796.txt";
test_data_files[2797] = "test_data_2797.txt";
test_data_files[2798] = "test_data_2798.txt";
test_data_files[2799] = "test_data_2799.txt";
test_data_files[2800] = "test_data_2800.txt";
test_data_files[2801] = "test_data_2801.txt";
test_data_files[2802] = "test_data_2802.txt";
test_data_files[2803] = "test_data_2803.txt";
test_data_files[2804] = "test_data_2804.txt";
test_data_files[2805] = "test_data_2805.txt";
test_data_files[2806] = "test_data_2806.txt";
test_data_files[2807] = "test_data_2807.txt";
test_data_files[2808] = "test_data_2808.txt";
test_data_files[2809] = "test_data_2809.txt";
test_data_files[2810] = "test_data_2810.txt";
test_data_files[2811] = "test_data_2811.txt";
test_data_files[2812] = "test_data_2812.txt";
test_data_files[2813] = "test_data_2813.txt";
test_data_files[2814] = "test_data_2814.txt";
test_data_files[2815] = "test_data_2815.txt";
test_data_files[2816] = "test_data_2816.txt";
test_data_files[2817] = "test_data_2817.txt";
test_data_files[2818] = "test_data_2818.txt";
test_data_files[2819] = "test_data_2819.txt";
test_data_files[2820] = "test_data_2820.txt";
test_data_files[2821] = "test_data_2821.txt";
test_data_files[2822] = "test_data_2822.txt";
test_data_files[2823] = "test_data_2823.txt";
test_data_files[2824] = "test_data_2824.txt";
test_data_files[2825] = "test_data_2825.txt";
test_data_files[2826] = "test_data_2826.txt";
test_data_files[2827] = "test_data_2827.txt";
test_data_files[2828] = "test_data_2828.txt";
test_data_files[2829] = "test_data_2829.txt";
test_data_files[2830] = "test_data_2830.txt";
test_data_files[2831] = "test_data_2831.txt";
test_data_files[2832] = "test_data_2832.txt";
test_data_files[2833] = "test_data_2833.txt";
test_data_files[2834] = "test_data_2834.txt";
test_data_files[2835] = "test_data_2835.txt";
test_data_files[2836] = "test_data_2836.txt";
test_data_files[2837] = "test_data_2837.txt";
test_data_files[2838] = "test_data_2838.txt";
test_data_files[2839] = "test_data_2839.txt";
test_data_files[2840] = "test_data_2840.txt";
test_data_files[2841] = "test_data_2841.txt";
test_data_files[2842] = "test_data_2842.txt";
test_data_files[2843] = "test_data_2843.txt";
test_data_files[2844] = "test_data_2844.txt";
test_data_files[2845] = "test_data_2845.txt";
test_data_files[2846] = "test_data_2846.txt";
test_data_files[2847] = "test_data_2847.txt";
test_data_files[2848] = "test_data_2848.txt";
test_data_files[2849] = "test_data_2849.txt";
test_data_files[2850] = "test_data_2850.txt";
test_data_files[2851] = "test_data_2851.txt";
test_data_files[2852] = "test_data_2852.txt";
test_data_files[2853] = "test_data_2853.txt";
test_data_files[2854] = "test_data_2854.txt";
test_data_files[2855] = "test_data_2855.txt";
test_data_files[2856] = "test_data_2856.txt";
test_data_files[2857] = "test_data_2857.txt";
test_data_files[2858] = "test_data_2858.txt";
test_data_files[2859] = "test_data_2859.txt";
test_data_files[2860] = "test_data_2860.txt";
test_data_files[2861] = "test_data_2861.txt";
test_data_files[2862] = "test_data_2862.txt";
test_data_files[2863] = "test_data_2863.txt";
test_data_files[2864] = "test_data_2864.txt";
test_data_files[2865] = "test_data_2865.txt";
test_data_files[2866] = "test_data_2866.txt";
test_data_files[2867] = "test_data_2867.txt";
test_data_files[2868] = "test_data_2868.txt";
test_data_files[2869] = "test_data_2869.txt";
test_data_files[2870] = "test_data_2870.txt";
test_data_files[2871] = "test_data_2871.txt";
test_data_files[2872] = "test_data_2872.txt";
test_data_files[2873] = "test_data_2873.txt";
test_data_files[2874] = "test_data_2874.txt";
test_data_files[2875] = "test_data_2875.txt";
test_data_files[2876] = "test_data_2876.txt";
test_data_files[2877] = "test_data_2877.txt";
test_data_files[2878] = "test_data_2878.txt";
test_data_files[2879] = "test_data_2879.txt";
test_data_files[2880] = "test_data_2880.txt";
test_data_files[2881] = "test_data_2881.txt";
test_data_files[2882] = "test_data_2882.txt";
test_data_files[2883] = "test_data_2883.txt";
test_data_files[2884] = "test_data_2884.txt";
test_data_files[2885] = "test_data_2885.txt";
test_data_files[2886] = "test_data_2886.txt";
test_data_files[2887] = "test_data_2887.txt";
test_data_files[2888] = "test_data_2888.txt";
test_data_files[2889] = "test_data_2889.txt";
test_data_files[2890] = "test_data_2890.txt";
test_data_files[2891] = "test_data_2891.txt";
test_data_files[2892] = "test_data_2892.txt";
test_data_files[2893] = "test_data_2893.txt";
test_data_files[2894] = "test_data_2894.txt";
test_data_files[2895] = "test_data_2895.txt";
test_data_files[2896] = "test_data_2896.txt";
test_data_files[2897] = "test_data_2897.txt";
test_data_files[2898] = "test_data_2898.txt";
test_data_files[2899] = "test_data_2899.txt";
test_data_files[2900] = "test_data_2900.txt";
test_data_files[2901] = "test_data_2901.txt";
test_data_files[2902] = "test_data_2902.txt";
test_data_files[2903] = "test_data_2903.txt";
test_data_files[2904] = "test_data_2904.txt";
test_data_files[2905] = "test_data_2905.txt";
test_data_files[2906] = "test_data_2906.txt";
test_data_files[2907] = "test_data_2907.txt";
test_data_files[2908] = "test_data_2908.txt";
test_data_files[2909] = "test_data_2909.txt";
test_data_files[2910] = "test_data_2910.txt";
test_data_files[2911] = "test_data_2911.txt";
test_data_files[2912] = "test_data_2912.txt";
test_data_files[2913] = "test_data_2913.txt";
test_data_files[2914] = "test_data_2914.txt";
test_data_files[2915] = "test_data_2915.txt";
test_data_files[2916] = "test_data_2916.txt";
test_data_files[2917] = "test_data_2917.txt";
test_data_files[2918] = "test_data_2918.txt";
test_data_files[2919] = "test_data_2919.txt";
test_data_files[2920] = "test_data_2920.txt";
test_data_files[2921] = "test_data_2921.txt";
test_data_files[2922] = "test_data_2922.txt";
test_data_files[2923] = "test_data_2923.txt";
test_data_files[2924] = "test_data_2924.txt";
test_data_files[2925] = "test_data_2925.txt";
test_data_files[2926] = "test_data_2926.txt";
test_data_files[2927] = "test_data_2927.txt";
test_data_files[2928] = "test_data_2928.txt";
test_data_files[2929] = "test_data_2929.txt";
test_data_files[2930] = "test_data_2930.txt";
test_data_files[2931] = "test_data_2931.txt";
test_data_files[2932] = "test_data_2932.txt";
test_data_files[2933] = "test_data_2933.txt";
test_data_files[2934] = "test_data_2934.txt";
test_data_files[2935] = "test_data_2935.txt";
test_data_files[2936] = "test_data_2936.txt";
test_data_files[2937] = "test_data_2937.txt";
test_data_files[2938] = "test_data_2938.txt";
test_data_files[2939] = "test_data_2939.txt";
test_data_files[2940] = "test_data_2940.txt";
test_data_files[2941] = "test_data_2941.txt";
test_data_files[2942] = "test_data_2942.txt";
test_data_files[2943] = "test_data_2943.txt";
test_data_files[2944] = "test_data_2944.txt";
test_data_files[2945] = "test_data_2945.txt";
test_data_files[2946] = "test_data_2946.txt";
test_data_files[2947] = "test_data_2947.txt";
test_data_files[2948] = "test_data_2948.txt";
test_data_files[2949] = "test_data_2949.txt";
test_data_files[2950] = "test_data_2950.txt";
test_data_files[2951] = "test_data_2951.txt";
test_data_files[2952] = "test_data_2952.txt";
test_data_files[2953] = "test_data_2953.txt";
test_data_files[2954] = "test_data_2954.txt";
test_data_files[2955] = "test_data_2955.txt";
test_data_files[2956] = "test_data_2956.txt";
test_data_files[2957] = "test_data_2957.txt";
test_data_files[2958] = "test_data_2958.txt";
test_data_files[2959] = "test_data_2959.txt";
test_data_files[2960] = "test_data_2960.txt";
test_data_files[2961] = "test_data_2961.txt";
test_data_files[2962] = "test_data_2962.txt";
test_data_files[2963] = "test_data_2963.txt";
test_data_files[2964] = "test_data_2964.txt";
test_data_files[2965] = "test_data_2965.txt";
test_data_files[2966] = "test_data_2966.txt";
test_data_files[2967] = "test_data_2967.txt";
test_data_files[2968] = "test_data_2968.txt";
test_data_files[2969] = "test_data_2969.txt";
test_data_files[2970] = "test_data_2970.txt";
test_data_files[2971] = "test_data_2971.txt";
test_data_files[2972] = "test_data_2972.txt";
test_data_files[2973] = "test_data_2973.txt";
test_data_files[2974] = "test_data_2974.txt";
test_data_files[2975] = "test_data_2975.txt";
test_data_files[2976] = "test_data_2976.txt";
test_data_files[2977] = "test_data_2977.txt";
test_data_files[2978] = "test_data_2978.txt";
test_data_files[2979] = "test_data_2979.txt";
test_data_files[2980] = "test_data_2980.txt";
test_data_files[2981] = "test_data_2981.txt";
test_data_files[2982] = "test_data_2982.txt";
test_data_files[2983] = "test_data_2983.txt";
test_data_files[2984] = "test_data_2984.txt";
test_data_files[2985] = "test_data_2985.txt";
test_data_files[2986] = "test_data_2986.txt";
test_data_files[2987] = "test_data_2987.txt";
test_data_files[2988] = "test_data_2988.txt";
test_data_files[2989] = "test_data_2989.txt";
test_data_files[2990] = "test_data_2990.txt";
test_data_files[2991] = "test_data_2991.txt";
test_data_files[2992] = "test_data_2992.txt";
test_data_files[2993] = "test_data_2993.txt";
test_data_files[2994] = "test_data_2994.txt";
test_data_files[2995] = "test_data_2995.txt";
test_data_files[2996] = "test_data_2996.txt";
test_data_files[2997] = "test_data_2997.txt";
test_data_files[2998] = "test_data_2998.txt";
test_data_files[2999] = "test_data_2999.txt";
test_data_files[3000] = "test_data_3000.txt";
test_data_files[3001] = "test_data_3001.txt";
test_data_files[3002] = "test_data_3002.txt";
test_data_files[3003] = "test_data_3003.txt";
test_data_files[3004] = "test_data_3004.txt";
test_data_files[3005] = "test_data_3005.txt";
test_data_files[3006] = "test_data_3006.txt";
test_data_files[3007] = "test_data_3007.txt";
test_data_files[3008] = "test_data_3008.txt";
test_data_files[3009] = "test_data_3009.txt";
test_data_files[3010] = "test_data_3010.txt";
test_data_files[3011] = "test_data_3011.txt";
test_data_files[3012] = "test_data_3012.txt";
test_data_files[3013] = "test_data_3013.txt";
test_data_files[3014] = "test_data_3014.txt";
test_data_files[3015] = "test_data_3015.txt";
test_data_files[3016] = "test_data_3016.txt";
test_data_files[3017] = "test_data_3017.txt";
test_data_files[3018] = "test_data_3018.txt";
test_data_files[3019] = "test_data_3019.txt";
test_data_files[3020] = "test_data_3020.txt";
test_data_files[3021] = "test_data_3021.txt";
test_data_files[3022] = "test_data_3022.txt";
test_data_files[3023] = "test_data_3023.txt";
test_data_files[3024] = "test_data_3024.txt";
test_data_files[3025] = "test_data_3025.txt";
test_data_files[3026] = "test_data_3026.txt";
test_data_files[3027] = "test_data_3027.txt";
test_data_files[3028] = "test_data_3028.txt";
test_data_files[3029] = "test_data_3029.txt";
test_data_files[3030] = "test_data_3030.txt";
test_data_files[3031] = "test_data_3031.txt";
test_data_files[3032] = "test_data_3032.txt";
test_data_files[3033] = "test_data_3033.txt";
test_data_files[3034] = "test_data_3034.txt";
test_data_files[3035] = "test_data_3035.txt";
test_data_files[3036] = "test_data_3036.txt";
test_data_files[3037] = "test_data_3037.txt";
test_data_files[3038] = "test_data_3038.txt";
test_data_files[3039] = "test_data_3039.txt";
test_data_files[3040] = "test_data_3040.txt";
test_data_files[3041] = "test_data_3041.txt";
test_data_files[3042] = "test_data_3042.txt";
test_data_files[3043] = "test_data_3043.txt";
test_data_files[3044] = "test_data_3044.txt";
test_data_files[3045] = "test_data_3045.txt";
test_data_files[3046] = "test_data_3046.txt";
test_data_files[3047] = "test_data_3047.txt";
test_data_files[3048] = "test_data_3048.txt";
test_data_files[3049] = "test_data_3049.txt";
test_data_files[3050] = "test_data_3050.txt";
test_data_files[3051] = "test_data_3051.txt";
test_data_files[3052] = "test_data_3052.txt";
test_data_files[3053] = "test_data_3053.txt";
test_data_files[3054] = "test_data_3054.txt";
test_data_files[3055] = "test_data_3055.txt";
test_data_files[3056] = "test_data_3056.txt";
test_data_files[3057] = "test_data_3057.txt";
test_data_files[3058] = "test_data_3058.txt";
test_data_files[3059] = "test_data_3059.txt";
test_data_files[3060] = "test_data_3060.txt";
test_data_files[3061] = "test_data_3061.txt";
test_data_files[3062] = "test_data_3062.txt";
test_data_files[3063] = "test_data_3063.txt";
test_data_files[3064] = "test_data_3064.txt";
test_data_files[3065] = "test_data_3065.txt";
test_data_files[3066] = "test_data_3066.txt";
test_data_files[3067] = "test_data_3067.txt";
test_data_files[3068] = "test_data_3068.txt";
test_data_files[3069] = "test_data_3069.txt";
test_data_files[3070] = "test_data_3070.txt";
test_data_files[3071] = "test_data_3071.txt";
test_data_files[3072] = "test_data_3072.txt";
test_data_files[3073] = "test_data_3073.txt";
test_data_files[3074] = "test_data_3074.txt";
test_data_files[3075] = "test_data_3075.txt";
test_data_files[3076] = "test_data_3076.txt";
test_data_files[3077] = "test_data_3077.txt";
test_data_files[3078] = "test_data_3078.txt";
test_data_files[3079] = "test_data_3079.txt";
test_data_files[3080] = "test_data_3080.txt";
test_data_files[3081] = "test_data_3081.txt";
test_data_files[3082] = "test_data_3082.txt";
test_data_files[3083] = "test_data_3083.txt";
test_data_files[3084] = "test_data_3084.txt";
test_data_files[3085] = "test_data_3085.txt";
test_data_files[3086] = "test_data_3086.txt";
test_data_files[3087] = "test_data_3087.txt";
test_data_files[3088] = "test_data_3088.txt";
test_data_files[3089] = "test_data_3089.txt";
test_data_files[3090] = "test_data_3090.txt";
test_data_files[3091] = "test_data_3091.txt";
test_data_files[3092] = "test_data_3092.txt";
test_data_files[3093] = "test_data_3093.txt";
test_data_files[3094] = "test_data_3094.txt";
test_data_files[3095] = "test_data_3095.txt";
test_data_files[3096] = "test_data_3096.txt";
test_data_files[3097] = "test_data_3097.txt";
test_data_files[3098] = "test_data_3098.txt";
test_data_files[3099] = "test_data_3099.txt";
test_data_files[3100] = "test_data_3100.txt";
test_data_files[3101] = "test_data_3101.txt";
test_data_files[3102] = "test_data_3102.txt";
test_data_files[3103] = "test_data_3103.txt";
test_data_files[3104] = "test_data_3104.txt";
test_data_files[3105] = "test_data_3105.txt";
test_data_files[3106] = "test_data_3106.txt";
test_data_files[3107] = "test_data_3107.txt";
test_data_files[3108] = "test_data_3108.txt";
test_data_files[3109] = "test_data_3109.txt";
test_data_files[3110] = "test_data_3110.txt";
test_data_files[3111] = "test_data_3111.txt";
test_data_files[3112] = "test_data_3112.txt";
test_data_files[3113] = "test_data_3113.txt";
test_data_files[3114] = "test_data_3114.txt";
test_data_files[3115] = "test_data_3115.txt";
test_data_files[3116] = "test_data_3116.txt";
test_data_files[3117] = "test_data_3117.txt";
test_data_files[3118] = "test_data_3118.txt";
test_data_files[3119] = "test_data_3119.txt";
test_data_files[3120] = "test_data_3120.txt";
test_data_files[3121] = "test_data_3121.txt";
test_data_files[3122] = "test_data_3122.txt";
test_data_files[3123] = "test_data_3123.txt";
test_data_files[3124] = "test_data_3124.txt";
test_data_files[3125] = "test_data_3125.txt";
test_data_files[3126] = "test_data_3126.txt";
test_data_files[3127] = "test_data_3127.txt";
test_data_files[3128] = "test_data_3128.txt";
test_data_files[3129] = "test_data_3129.txt";
test_data_files[3130] = "test_data_3130.txt";
test_data_files[3131] = "test_data_3131.txt";
test_data_files[3132] = "test_data_3132.txt";
test_data_files[3133] = "test_data_3133.txt";
test_data_files[3134] = "test_data_3134.txt";
test_data_files[3135] = "test_data_3135.txt";
test_data_files[3136] = "test_data_3136.txt";
test_data_files[3137] = "test_data_3137.txt";
test_data_files[3138] = "test_data_3138.txt";
test_data_files[3139] = "test_data_3139.txt";
test_data_files[3140] = "test_data_3140.txt";
test_data_files[3141] = "test_data_3141.txt";
test_data_files[3142] = "test_data_3142.txt";
test_data_files[3143] = "test_data_3143.txt";
test_data_files[3144] = "test_data_3144.txt";
test_data_files[3145] = "test_data_3145.txt";
test_data_files[3146] = "test_data_3146.txt";
test_data_files[3147] = "test_data_3147.txt";
test_data_files[3148] = "test_data_3148.txt";
test_data_files[3149] = "test_data_3149.txt";
test_data_files[3150] = "test_data_3150.txt";
test_data_files[3151] = "test_data_3151.txt";
test_data_files[3152] = "test_data_3152.txt";
test_data_files[3153] = "test_data_3153.txt";
test_data_files[3154] = "test_data_3154.txt";
test_data_files[3155] = "test_data_3155.txt";
test_data_files[3156] = "test_data_3156.txt";
test_data_files[3157] = "test_data_3157.txt";
test_data_files[3158] = "test_data_3158.txt";
test_data_files[3159] = "test_data_3159.txt";
test_data_files[3160] = "test_data_3160.txt";
test_data_files[3161] = "test_data_3161.txt";
test_data_files[3162] = "test_data_3162.txt";
test_data_files[3163] = "test_data_3163.txt";
test_data_files[3164] = "test_data_3164.txt";
test_data_files[3165] = "test_data_3165.txt";
test_data_files[3166] = "test_data_3166.txt";
test_data_files[3167] = "test_data_3167.txt";
test_data_files[3168] = "test_data_3168.txt";
test_data_files[3169] = "test_data_3169.txt";
test_data_files[3170] = "test_data_3170.txt";
test_data_files[3171] = "test_data_3171.txt";
test_data_files[3172] = "test_data_3172.txt";
test_data_files[3173] = "test_data_3173.txt";
test_data_files[3174] = "test_data_3174.txt";
test_data_files[3175] = "test_data_3175.txt";
test_data_files[3176] = "test_data_3176.txt";
test_data_files[3177] = "test_data_3177.txt";
test_data_files[3178] = "test_data_3178.txt";
test_data_files[3179] = "test_data_3179.txt";
test_data_files[3180] = "test_data_3180.txt";
test_data_files[3181] = "test_data_3181.txt";
test_data_files[3182] = "test_data_3182.txt";
test_data_files[3183] = "test_data_3183.txt";
test_data_files[3184] = "test_data_3184.txt";
test_data_files[3185] = "test_data_3185.txt";
test_data_files[3186] = "test_data_3186.txt";
test_data_files[3187] = "test_data_3187.txt";
test_data_files[3188] = "test_data_3188.txt";
test_data_files[3189] = "test_data_3189.txt";
test_data_files[3190] = "test_data_3190.txt";
test_data_files[3191] = "test_data_3191.txt";
test_data_files[3192] = "test_data_3192.txt";
test_data_files[3193] = "test_data_3193.txt";
test_data_files[3194] = "test_data_3194.txt";
test_data_files[3195] = "test_data_3195.txt";
test_data_files[3196] = "test_data_3196.txt";
test_data_files[3197] = "test_data_3197.txt";
test_data_files[3198] = "test_data_3198.txt";
test_data_files[3199] = "test_data_3199.txt";
test_data_files[3200] = "test_data_3200.txt";
test_data_files[3201] = "test_data_3201.txt";
test_data_files[3202] = "test_data_3202.txt";
test_data_files[3203] = "test_data_3203.txt";
test_data_files[3204] = "test_data_3204.txt";
test_data_files[3205] = "test_data_3205.txt";
test_data_files[3206] = "test_data_3206.txt";
test_data_files[3207] = "test_data_3207.txt";
test_data_files[3208] = "test_data_3208.txt";
test_data_files[3209] = "test_data_3209.txt";
test_data_files[3210] = "test_data_3210.txt";
test_data_files[3211] = "test_data_3211.txt";
test_data_files[3212] = "test_data_3212.txt";
test_data_files[3213] = "test_data_3213.txt";
test_data_files[3214] = "test_data_3214.txt";
test_data_files[3215] = "test_data_3215.txt";
test_data_files[3216] = "test_data_3216.txt";
test_data_files[3217] = "test_data_3217.txt";
test_data_files[3218] = "test_data_3218.txt";
test_data_files[3219] = "test_data_3219.txt";
test_data_files[3220] = "test_data_3220.txt";
test_data_files[3221] = "test_data_3221.txt";
test_data_files[3222] = "test_data_3222.txt";
test_data_files[3223] = "test_data_3223.txt";
test_data_files[3224] = "test_data_3224.txt";
test_data_files[3225] = "test_data_3225.txt";
test_data_files[3226] = "test_data_3226.txt";
test_data_files[3227] = "test_data_3227.txt";
test_data_files[3228] = "test_data_3228.txt";
test_data_files[3229] = "test_data_3229.txt";
test_data_files[3230] = "test_data_3230.txt";
test_data_files[3231] = "test_data_3231.txt";
test_data_files[3232] = "test_data_3232.txt";
test_data_files[3233] = "test_data_3233.txt";
test_data_files[3234] = "test_data_3234.txt";
test_data_files[3235] = "test_data_3235.txt";
test_data_files[3236] = "test_data_3236.txt";
test_data_files[3237] = "test_data_3237.txt";
test_data_files[3238] = "test_data_3238.txt";
test_data_files[3239] = "test_data_3239.txt";
test_data_files[3240] = "test_data_3240.txt";
test_data_files[3241] = "test_data_3241.txt";
test_data_files[3242] = "test_data_3242.txt";
test_data_files[3243] = "test_data_3243.txt";
test_data_files[3244] = "test_data_3244.txt";
test_data_files[3245] = "test_data_3245.txt";
test_data_files[3246] = "test_data_3246.txt";
test_data_files[3247] = "test_data_3247.txt";
test_data_files[3248] = "test_data_3248.txt";
test_data_files[3249] = "test_data_3249.txt";
test_data_files[3250] = "test_data_3250.txt";
test_data_files[3251] = "test_data_3251.txt";
test_data_files[3252] = "test_data_3252.txt";
test_data_files[3253] = "test_data_3253.txt";
test_data_files[3254] = "test_data_3254.txt";
test_data_files[3255] = "test_data_3255.txt";
test_data_files[3256] = "test_data_3256.txt";
test_data_files[3257] = "test_data_3257.txt";
test_data_files[3258] = "test_data_3258.txt";
test_data_files[3259] = "test_data_3259.txt";
test_data_files[3260] = "test_data_3260.txt";
test_data_files[3261] = "test_data_3261.txt";
test_data_files[3262] = "test_data_3262.txt";
test_data_files[3263] = "test_data_3263.txt";
test_data_files[3264] = "test_data_3264.txt";
test_data_files[3265] = "test_data_3265.txt";
test_data_files[3266] = "test_data_3266.txt";
test_data_files[3267] = "test_data_3267.txt";
test_data_files[3268] = "test_data_3268.txt";
test_data_files[3269] = "test_data_3269.txt";
test_data_files[3270] = "test_data_3270.txt";
test_data_files[3271] = "test_data_3271.txt";
test_data_files[3272] = "test_data_3272.txt";
test_data_files[3273] = "test_data_3273.txt";
test_data_files[3274] = "test_data_3274.txt";
test_data_files[3275] = "test_data_3275.txt";
test_data_files[3276] = "test_data_3276.txt";
test_data_files[3277] = "test_data_3277.txt";
test_data_files[3278] = "test_data_3278.txt";
test_data_files[3279] = "test_data_3279.txt";
test_data_files[3280] = "test_data_3280.txt";
test_data_files[3281] = "test_data_3281.txt";
test_data_files[3282] = "test_data_3282.txt";
test_data_files[3283] = "test_data_3283.txt";
test_data_files[3284] = "test_data_3284.txt";
test_data_files[3285] = "test_data_3285.txt";
test_data_files[3286] = "test_data_3286.txt";
test_data_files[3287] = "test_data_3287.txt";
test_data_files[3288] = "test_data_3288.txt";
test_data_files[3289] = "test_data_3289.txt";
test_data_files[3290] = "test_data_3290.txt";
test_data_files[3291] = "test_data_3291.txt";
test_data_files[3292] = "test_data_3292.txt";
test_data_files[3293] = "test_data_3293.txt";
test_data_files[3294] = "test_data_3294.txt";
test_data_files[3295] = "test_data_3295.txt";
test_data_files[3296] = "test_data_3296.txt";
test_data_files[3297] = "test_data_3297.txt";
test_data_files[3298] = "test_data_3298.txt";
test_data_files[3299] = "test_data_3299.txt";
test_data_files[3300] = "test_data_3300.txt";
test_data_files[3301] = "test_data_3301.txt";
test_data_files[3302] = "test_data_3302.txt";
test_data_files[3303] = "test_data_3303.txt";
test_data_files[3304] = "test_data_3304.txt";
test_data_files[3305] = "test_data_3305.txt";
test_data_files[3306] = "test_data_3306.txt";
test_data_files[3307] = "test_data_3307.txt";
test_data_files[3308] = "test_data_3308.txt";
test_data_files[3309] = "test_data_3309.txt";
test_data_files[3310] = "test_data_3310.txt";
test_data_files[3311] = "test_data_3311.txt";
test_data_files[3312] = "test_data_3312.txt";
test_data_files[3313] = "test_data_3313.txt";
test_data_files[3314] = "test_data_3314.txt";
test_data_files[3315] = "test_data_3315.txt";
test_data_files[3316] = "test_data_3316.txt";
test_data_files[3317] = "test_data_3317.txt";
test_data_files[3318] = "test_data_3318.txt";
test_data_files[3319] = "test_data_3319.txt";
test_data_files[3320] = "test_data_3320.txt";
test_data_files[3321] = "test_data_3321.txt";
test_data_files[3322] = "test_data_3322.txt";
test_data_files[3323] = "test_data_3323.txt";
test_data_files[3324] = "test_data_3324.txt";
test_data_files[3325] = "test_data_3325.txt";
test_data_files[3326] = "test_data_3326.txt";
test_data_files[3327] = "test_data_3327.txt";
test_data_files[3328] = "test_data_3328.txt";
test_data_files[3329] = "test_data_3329.txt";
test_data_files[3330] = "test_data_3330.txt";
test_data_files[3331] = "test_data_3331.txt";
test_data_files[3332] = "test_data_3332.txt";
test_data_files[3333] = "test_data_3333.txt";
test_data_files[3334] = "test_data_3334.txt";
test_data_files[3335] = "test_data_3335.txt";
test_data_files[3336] = "test_data_3336.txt";
test_data_files[3337] = "test_data_3337.txt";
test_data_files[3338] = "test_data_3338.txt";
test_data_files[3339] = "test_data_3339.txt";
test_data_files[3340] = "test_data_3340.txt";
test_data_files[3341] = "test_data_3341.txt";
test_data_files[3342] = "test_data_3342.txt";
test_data_files[3343] = "test_data_3343.txt";
test_data_files[3344] = "test_data_3344.txt";
test_data_files[3345] = "test_data_3345.txt";
test_data_files[3346] = "test_data_3346.txt";
test_data_files[3347] = "test_data_3347.txt";
test_data_files[3348] = "test_data_3348.txt";
test_data_files[3349] = "test_data_3349.txt";
test_data_files[3350] = "test_data_3350.txt";
test_data_files[3351] = "test_data_3351.txt";
test_data_files[3352] = "test_data_3352.txt";
test_data_files[3353] = "test_data_3353.txt";
test_data_files[3354] = "test_data_3354.txt";
test_data_files[3355] = "test_data_3355.txt";
test_data_files[3356] = "test_data_3356.txt";
test_data_files[3357] = "test_data_3357.txt";
test_data_files[3358] = "test_data_3358.txt";
test_data_files[3359] = "test_data_3359.txt";
test_data_files[3360] = "test_data_3360.txt";
test_data_files[3361] = "test_data_3361.txt";
test_data_files[3362] = "test_data_3362.txt";
test_data_files[3363] = "test_data_3363.txt";
test_data_files[3364] = "test_data_3364.txt";
test_data_files[3365] = "test_data_3365.txt";
test_data_files[3366] = "test_data_3366.txt";
test_data_files[3367] = "test_data_3367.txt";
test_data_files[3368] = "test_data_3368.txt";
test_data_files[3369] = "test_data_3369.txt";
test_data_files[3370] = "test_data_3370.txt";
test_data_files[3371] = "test_data_3371.txt";
test_data_files[3372] = "test_data_3372.txt";
test_data_files[3373] = "test_data_3373.txt";
test_data_files[3374] = "test_data_3374.txt";
test_data_files[3375] = "test_data_3375.txt";
test_data_files[3376] = "test_data_3376.txt";
test_data_files[3377] = "test_data_3377.txt";
test_data_files[3378] = "test_data_3378.txt";
test_data_files[3379] = "test_data_3379.txt";
test_data_files[3380] = "test_data_3380.txt";
test_data_files[3381] = "test_data_3381.txt";
test_data_files[3382] = "test_data_3382.txt";
test_data_files[3383] = "test_data_3383.txt";
test_data_files[3384] = "test_data_3384.txt";
test_data_files[3385] = "test_data_3385.txt";
test_data_files[3386] = "test_data_3386.txt";
test_data_files[3387] = "test_data_3387.txt";
test_data_files[3388] = "test_data_3388.txt";
test_data_files[3389] = "test_data_3389.txt";
test_data_files[3390] = "test_data_3390.txt";
test_data_files[3391] = "test_data_3391.txt";
test_data_files[3392] = "test_data_3392.txt";
test_data_files[3393] = "test_data_3393.txt";
test_data_files[3394] = "test_data_3394.txt";
test_data_files[3395] = "test_data_3395.txt";
test_data_files[3396] = "test_data_3396.txt";
test_data_files[3397] = "test_data_3397.txt";
test_data_files[3398] = "test_data_3398.txt";
test_data_files[3399] = "test_data_3399.txt";
test_data_files[3400] = "test_data_3400.txt";
test_data_files[3401] = "test_data_3401.txt";
test_data_files[3402] = "test_data_3402.txt";
test_data_files[3403] = "test_data_3403.txt";
test_data_files[3404] = "test_data_3404.txt";
test_data_files[3405] = "test_data_3405.txt";
test_data_files[3406] = "test_data_3406.txt";
test_data_files[3407] = "test_data_3407.txt";
test_data_files[3408] = "test_data_3408.txt";
test_data_files[3409] = "test_data_3409.txt";
test_data_files[3410] = "test_data_3410.txt";
test_data_files[3411] = "test_data_3411.txt";
test_data_files[3412] = "test_data_3412.txt";
test_data_files[3413] = "test_data_3413.txt";
test_data_files[3414] = "test_data_3414.txt";
test_data_files[3415] = "test_data_3415.txt";
test_data_files[3416] = "test_data_3416.txt";
test_data_files[3417] = "test_data_3417.txt";
test_data_files[3418] = "test_data_3418.txt";
test_data_files[3419] = "test_data_3419.txt";
test_data_files[3420] = "test_data_3420.txt";
test_data_files[3421] = "test_data_3421.txt";
test_data_files[3422] = "test_data_3422.txt";
test_data_files[3423] = "test_data_3423.txt";
test_data_files[3424] = "test_data_3424.txt";
test_data_files[3425] = "test_data_3425.txt";
test_data_files[3426] = "test_data_3426.txt";
test_data_files[3427] = "test_data_3427.txt";
test_data_files[3428] = "test_data_3428.txt";
test_data_files[3429] = "test_data_3429.txt";
test_data_files[3430] = "test_data_3430.txt";
test_data_files[3431] = "test_data_3431.txt";
test_data_files[3432] = "test_data_3432.txt";
test_data_files[3433] = "test_data_3433.txt";
test_data_files[3434] = "test_data_3434.txt";
test_data_files[3435] = "test_data_3435.txt";
test_data_files[3436] = "test_data_3436.txt";
test_data_files[3437] = "test_data_3437.txt";
test_data_files[3438] = "test_data_3438.txt";
test_data_files[3439] = "test_data_3439.txt";
test_data_files[3440] = "test_data_3440.txt";
test_data_files[3441] = "test_data_3441.txt";
test_data_files[3442] = "test_data_3442.txt";
test_data_files[3443] = "test_data_3443.txt";
test_data_files[3444] = "test_data_3444.txt";
test_data_files[3445] = "test_data_3445.txt";
test_data_files[3446] = "test_data_3446.txt";
test_data_files[3447] = "test_data_3447.txt";
test_data_files[3448] = "test_data_3448.txt";
test_data_files[3449] = "test_data_3449.txt";
test_data_files[3450] = "test_data_3450.txt";
test_data_files[3451] = "test_data_3451.txt";
test_data_files[3452] = "test_data_3452.txt";
test_data_files[3453] = "test_data_3453.txt";
test_data_files[3454] = "test_data_3454.txt";
test_data_files[3455] = "test_data_3455.txt";
test_data_files[3456] = "test_data_3456.txt";
test_data_files[3457] = "test_data_3457.txt";
test_data_files[3458] = "test_data_3458.txt";
test_data_files[3459] = "test_data_3459.txt";
test_data_files[3460] = "test_data_3460.txt";
test_data_files[3461] = "test_data_3461.txt";
test_data_files[3462] = "test_data_3462.txt";
test_data_files[3463] = "test_data_3463.txt";
test_data_files[3464] = "test_data_3464.txt";
test_data_files[3465] = "test_data_3465.txt";
test_data_files[3466] = "test_data_3466.txt";
test_data_files[3467] = "test_data_3467.txt";
test_data_files[3468] = "test_data_3468.txt";
test_data_files[3469] = "test_data_3469.txt";
test_data_files[3470] = "test_data_3470.txt";
test_data_files[3471] = "test_data_3471.txt";
test_data_files[3472] = "test_data_3472.txt";
test_data_files[3473] = "test_data_3473.txt";
test_data_files[3474] = "test_data_3474.txt";
test_data_files[3475] = "test_data_3475.txt";
test_data_files[3476] = "test_data_3476.txt";
test_data_files[3477] = "test_data_3477.txt";
test_data_files[3478] = "test_data_3478.txt";
test_data_files[3479] = "test_data_3479.txt";
test_data_files[3480] = "test_data_3480.txt";
test_data_files[3481] = "test_data_3481.txt";
test_data_files[3482] = "test_data_3482.txt";
test_data_files[3483] = "test_data_3483.txt";
test_data_files[3484] = "test_data_3484.txt";
test_data_files[3485] = "test_data_3485.txt";
test_data_files[3486] = "test_data_3486.txt";
test_data_files[3487] = "test_data_3487.txt";
test_data_files[3488] = "test_data_3488.txt";
test_data_files[3489] = "test_data_3489.txt";
test_data_files[3490] = "test_data_3490.txt";
test_data_files[3491] = "test_data_3491.txt";
test_data_files[3492] = "test_data_3492.txt";
test_data_files[3493] = "test_data_3493.txt";
test_data_files[3494] = "test_data_3494.txt";
test_data_files[3495] = "test_data_3495.txt";
test_data_files[3496] = "test_data_3496.txt";
test_data_files[3497] = "test_data_3497.txt";
test_data_files[3498] = "test_data_3498.txt";
test_data_files[3499] = "test_data_3499.txt";
test_data_files[3500] = "test_data_3500.txt";
test_data_files[3501] = "test_data_3501.txt";
test_data_files[3502] = "test_data_3502.txt";
test_data_files[3503] = "test_data_3503.txt";
test_data_files[3504] = "test_data_3504.txt";
test_data_files[3505] = "test_data_3505.txt";
test_data_files[3506] = "test_data_3506.txt";
test_data_files[3507] = "test_data_3507.txt";
test_data_files[3508] = "test_data_3508.txt";
test_data_files[3509] = "test_data_3509.txt";
test_data_files[3510] = "test_data_3510.txt";
test_data_files[3511] = "test_data_3511.txt";
test_data_files[3512] = "test_data_3512.txt";
test_data_files[3513] = "test_data_3513.txt";
test_data_files[3514] = "test_data_3514.txt";
test_data_files[3515] = "test_data_3515.txt";
test_data_files[3516] = "test_data_3516.txt";
test_data_files[3517] = "test_data_3517.txt";
test_data_files[3518] = "test_data_3518.txt";
test_data_files[3519] = "test_data_3519.txt";
test_data_files[3520] = "test_data_3520.txt";
test_data_files[3521] = "test_data_3521.txt";
test_data_files[3522] = "test_data_3522.txt";
test_data_files[3523] = "test_data_3523.txt";
test_data_files[3524] = "test_data_3524.txt";
test_data_files[3525] = "test_data_3525.txt";
test_data_files[3526] = "test_data_3526.txt";
test_data_files[3527] = "test_data_3527.txt";
test_data_files[3528] = "test_data_3528.txt";
test_data_files[3529] = "test_data_3529.txt";
test_data_files[3530] = "test_data_3530.txt";
test_data_files[3531] = "test_data_3531.txt";
test_data_files[3532] = "test_data_3532.txt";
test_data_files[3533] = "test_data_3533.txt";
test_data_files[3534] = "test_data_3534.txt";
test_data_files[3535] = "test_data_3535.txt";
test_data_files[3536] = "test_data_3536.txt";
test_data_files[3537] = "test_data_3537.txt";
test_data_files[3538] = "test_data_3538.txt";
test_data_files[3539] = "test_data_3539.txt";
test_data_files[3540] = "test_data_3540.txt";
test_data_files[3541] = "test_data_3541.txt";
test_data_files[3542] = "test_data_3542.txt";
test_data_files[3543] = "test_data_3543.txt";
test_data_files[3544] = "test_data_3544.txt";
test_data_files[3545] = "test_data_3545.txt";
test_data_files[3546] = "test_data_3546.txt";
test_data_files[3547] = "test_data_3547.txt";
test_data_files[3548] = "test_data_3548.txt";
test_data_files[3549] = "test_data_3549.txt";
test_data_files[3550] = "test_data_3550.txt";
test_data_files[3551] = "test_data_3551.txt";
test_data_files[3552] = "test_data_3552.txt";
test_data_files[3553] = "test_data_3553.txt";
test_data_files[3554] = "test_data_3554.txt";
test_data_files[3555] = "test_data_3555.txt";
test_data_files[3556] = "test_data_3556.txt";
test_data_files[3557] = "test_data_3557.txt";
test_data_files[3558] = "test_data_3558.txt";
test_data_files[3559] = "test_data_3559.txt";
test_data_files[3560] = "test_data_3560.txt";
test_data_files[3561] = "test_data_3561.txt";
test_data_files[3562] = "test_data_3562.txt";
test_data_files[3563] = "test_data_3563.txt";
test_data_files[3564] = "test_data_3564.txt";
test_data_files[3565] = "test_data_3565.txt";
test_data_files[3566] = "test_data_3566.txt";
test_data_files[3567] = "test_data_3567.txt";
test_data_files[3568] = "test_data_3568.txt";
test_data_files[3569] = "test_data_3569.txt";
test_data_files[3570] = "test_data_3570.txt";
test_data_files[3571] = "test_data_3571.txt";
test_data_files[3572] = "test_data_3572.txt";
test_data_files[3573] = "test_data_3573.txt";
test_data_files[3574] = "test_data_3574.txt";
test_data_files[3575] = "test_data_3575.txt";
test_data_files[3576] = "test_data_3576.txt";
test_data_files[3577] = "test_data_3577.txt";
test_data_files[3578] = "test_data_3578.txt";
test_data_files[3579] = "test_data_3579.txt";
test_data_files[3580] = "test_data_3580.txt";
test_data_files[3581] = "test_data_3581.txt";
test_data_files[3582] = "test_data_3582.txt";
test_data_files[3583] = "test_data_3583.txt";
test_data_files[3584] = "test_data_3584.txt";
test_data_files[3585] = "test_data_3585.txt";
test_data_files[3586] = "test_data_3586.txt";
test_data_files[3587] = "test_data_3587.txt";
test_data_files[3588] = "test_data_3588.txt";
test_data_files[3589] = "test_data_3589.txt";
test_data_files[3590] = "test_data_3590.txt";
test_data_files[3591] = "test_data_3591.txt";
test_data_files[3592] = "test_data_3592.txt";
test_data_files[3593] = "test_data_3593.txt";
test_data_files[3594] = "test_data_3594.txt";
test_data_files[3595] = "test_data_3595.txt";
test_data_files[3596] = "test_data_3596.txt";
test_data_files[3597] = "test_data_3597.txt";
test_data_files[3598] = "test_data_3598.txt";
test_data_files[3599] = "test_data_3599.txt";
test_data_files[3600] = "test_data_3600.txt";
test_data_files[3601] = "test_data_3601.txt";
test_data_files[3602] = "test_data_3602.txt";
test_data_files[3603] = "test_data_3603.txt";
test_data_files[3604] = "test_data_3604.txt";
test_data_files[3605] = "test_data_3605.txt";
test_data_files[3606] = "test_data_3606.txt";
test_data_files[3607] = "test_data_3607.txt";
test_data_files[3608] = "test_data_3608.txt";
test_data_files[3609] = "test_data_3609.txt";
test_data_files[3610] = "test_data_3610.txt";
test_data_files[3611] = "test_data_3611.txt";
test_data_files[3612] = "test_data_3612.txt";
test_data_files[3613] = "test_data_3613.txt";
test_data_files[3614] = "test_data_3614.txt";
test_data_files[3615] = "test_data_3615.txt";
test_data_files[3616] = "test_data_3616.txt";
test_data_files[3617] = "test_data_3617.txt";
test_data_files[3618] = "test_data_3618.txt";
test_data_files[3619] = "test_data_3619.txt";
test_data_files[3620] = "test_data_3620.txt";
test_data_files[3621] = "test_data_3621.txt";
test_data_files[3622] = "test_data_3622.txt";
test_data_files[3623] = "test_data_3623.txt";
test_data_files[3624] = "test_data_3624.txt";
test_data_files[3625] = "test_data_3625.txt";
test_data_files[3626] = "test_data_3626.txt";
test_data_files[3627] = "test_data_3627.txt";
test_data_files[3628] = "test_data_3628.txt";
test_data_files[3629] = "test_data_3629.txt";
test_data_files[3630] = "test_data_3630.txt";
test_data_files[3631] = "test_data_3631.txt";
test_data_files[3632] = "test_data_3632.txt";
test_data_files[3633] = "test_data_3633.txt";
test_data_files[3634] = "test_data_3634.txt";
test_data_files[3635] = "test_data_3635.txt";
test_data_files[3636] = "test_data_3636.txt";
test_data_files[3637] = "test_data_3637.txt";
test_data_files[3638] = "test_data_3638.txt";
test_data_files[3639] = "test_data_3639.txt";
test_data_files[3640] = "test_data_3640.txt";
test_data_files[3641] = "test_data_3641.txt";
test_data_files[3642] = "test_data_3642.txt";
test_data_files[3643] = "test_data_3643.txt";
test_data_files[3644] = "test_data_3644.txt";
test_data_files[3645] = "test_data_3645.txt";
test_data_files[3646] = "test_data_3646.txt";
test_data_files[3647] = "test_data_3647.txt";
test_data_files[3648] = "test_data_3648.txt";
test_data_files[3649] = "test_data_3649.txt";
test_data_files[3650] = "test_data_3650.txt";
test_data_files[3651] = "test_data_3651.txt";
test_data_files[3652] = "test_data_3652.txt";
test_data_files[3653] = "test_data_3653.txt";
test_data_files[3654] = "test_data_3654.txt";
test_data_files[3655] = "test_data_3655.txt";
test_data_files[3656] = "test_data_3656.txt";
test_data_files[3657] = "test_data_3657.txt";
test_data_files[3658] = "test_data_3658.txt";
test_data_files[3659] = "test_data_3659.txt";
test_data_files[3660] = "test_data_3660.txt";
test_data_files[3661] = "test_data_3661.txt";
test_data_files[3662] = "test_data_3662.txt";
test_data_files[3663] = "test_data_3663.txt";
test_data_files[3664] = "test_data_3664.txt";
test_data_files[3665] = "test_data_3665.txt";
test_data_files[3666] = "test_data_3666.txt";
test_data_files[3667] = "test_data_3667.txt";
test_data_files[3668] = "test_data_3668.txt";
test_data_files[3669] = "test_data_3669.txt";
test_data_files[3670] = "test_data_3670.txt";
test_data_files[3671] = "test_data_3671.txt";
test_data_files[3672] = "test_data_3672.txt";
test_data_files[3673] = "test_data_3673.txt";
test_data_files[3674] = "test_data_3674.txt";
test_data_files[3675] = "test_data_3675.txt";
test_data_files[3676] = "test_data_3676.txt";
test_data_files[3677] = "test_data_3677.txt";
test_data_files[3678] = "test_data_3678.txt";
test_data_files[3679] = "test_data_3679.txt";
test_data_files[3680] = "test_data_3680.txt";
test_data_files[3681] = "test_data_3681.txt";
test_data_files[3682] = "test_data_3682.txt";
test_data_files[3683] = "test_data_3683.txt";
test_data_files[3684] = "test_data_3684.txt";
test_data_files[3685] = "test_data_3685.txt";
test_data_files[3686] = "test_data_3686.txt";
test_data_files[3687] = "test_data_3687.txt";
test_data_files[3688] = "test_data_3688.txt";
test_data_files[3689] = "test_data_3689.txt";
test_data_files[3690] = "test_data_3690.txt";
test_data_files[3691] = "test_data_3691.txt";
test_data_files[3692] = "test_data_3692.txt";
test_data_files[3693] = "test_data_3693.txt";
test_data_files[3694] = "test_data_3694.txt";
test_data_files[3695] = "test_data_3695.txt";
test_data_files[3696] = "test_data_3696.txt";
test_data_files[3697] = "test_data_3697.txt";
test_data_files[3698] = "test_data_3698.txt";
test_data_files[3699] = "test_data_3699.txt";
test_data_files[3700] = "test_data_3700.txt";
test_data_files[3701] = "test_data_3701.txt";
test_data_files[3702] = "test_data_3702.txt";
test_data_files[3703] = "test_data_3703.txt";
test_data_files[3704] = "test_data_3704.txt";
test_data_files[3705] = "test_data_3705.txt";
test_data_files[3706] = "test_data_3706.txt";
test_data_files[3707] = "test_data_3707.txt";
test_data_files[3708] = "test_data_3708.txt";
test_data_files[3709] = "test_data_3709.txt";
test_data_files[3710] = "test_data_3710.txt";
test_data_files[3711] = "test_data_3711.txt";
test_data_files[3712] = "test_data_3712.txt";
test_data_files[3713] = "test_data_3713.txt";
test_data_files[3714] = "test_data_3714.txt";
test_data_files[3715] = "test_data_3715.txt";
test_data_files[3716] = "test_data_3716.txt";
test_data_files[3717] = "test_data_3717.txt";
test_data_files[3718] = "test_data_3718.txt";
test_data_files[3719] = "test_data_3719.txt";
test_data_files[3720] = "test_data_3720.txt";
test_data_files[3721] = "test_data_3721.txt";
test_data_files[3722] = "test_data_3722.txt";
test_data_files[3723] = "test_data_3723.txt";
test_data_files[3724] = "test_data_3724.txt";
test_data_files[3725] = "test_data_3725.txt";
test_data_files[3726] = "test_data_3726.txt";
test_data_files[3727] = "test_data_3727.txt";
test_data_files[3728] = "test_data_3728.txt";
test_data_files[3729] = "test_data_3729.txt";
test_data_files[3730] = "test_data_3730.txt";
test_data_files[3731] = "test_data_3731.txt";
test_data_files[3732] = "test_data_3732.txt";
test_data_files[3733] = "test_data_3733.txt";
test_data_files[3734] = "test_data_3734.txt";
test_data_files[3735] = "test_data_3735.txt";
test_data_files[3736] = "test_data_3736.txt";
test_data_files[3737] = "test_data_3737.txt";
test_data_files[3738] = "test_data_3738.txt";
test_data_files[3739] = "test_data_3739.txt";
test_data_files[3740] = "test_data_3740.txt";
test_data_files[3741] = "test_data_3741.txt";
test_data_files[3742] = "test_data_3742.txt";
test_data_files[3743] = "test_data_3743.txt";
test_data_files[3744] = "test_data_3744.txt";
test_data_files[3745] = "test_data_3745.txt";
test_data_files[3746] = "test_data_3746.txt";
test_data_files[3747] = "test_data_3747.txt";
test_data_files[3748] = "test_data_3748.txt";
test_data_files[3749] = "test_data_3749.txt";
test_data_files[3750] = "test_data_3750.txt";
test_data_files[3751] = "test_data_3751.txt";
test_data_files[3752] = "test_data_3752.txt";
test_data_files[3753] = "test_data_3753.txt";
test_data_files[3754] = "test_data_3754.txt";
test_data_files[3755] = "test_data_3755.txt";
test_data_files[3756] = "test_data_3756.txt";
test_data_files[3757] = "test_data_3757.txt";
test_data_files[3758] = "test_data_3758.txt";
test_data_files[3759] = "test_data_3759.txt";
test_data_files[3760] = "test_data_3760.txt";
test_data_files[3761] = "test_data_3761.txt";
test_data_files[3762] = "test_data_3762.txt";
test_data_files[3763] = "test_data_3763.txt";
test_data_files[3764] = "test_data_3764.txt";
test_data_files[3765] = "test_data_3765.txt";
test_data_files[3766] = "test_data_3766.txt";
test_data_files[3767] = "test_data_3767.txt";
test_data_files[3768] = "test_data_3768.txt";
test_data_files[3769] = "test_data_3769.txt";
test_data_files[3770] = "test_data_3770.txt";
test_data_files[3771] = "test_data_3771.txt";
test_data_files[3772] = "test_data_3772.txt";
test_data_files[3773] = "test_data_3773.txt";
test_data_files[3774] = "test_data_3774.txt";
test_data_files[3775] = "test_data_3775.txt";
test_data_files[3776] = "test_data_3776.txt";
test_data_files[3777] = "test_data_3777.txt";
test_data_files[3778] = "test_data_3778.txt";
test_data_files[3779] = "test_data_3779.txt";
test_data_files[3780] = "test_data_3780.txt";
test_data_files[3781] = "test_data_3781.txt";
test_data_files[3782] = "test_data_3782.txt";
test_data_files[3783] = "test_data_3783.txt";
test_data_files[3784] = "test_data_3784.txt";
test_data_files[3785] = "test_data_3785.txt";
test_data_files[3786] = "test_data_3786.txt";
test_data_files[3787] = "test_data_3787.txt";
test_data_files[3788] = "test_data_3788.txt";
test_data_files[3789] = "test_data_3789.txt";
test_data_files[3790] = "test_data_3790.txt";
test_data_files[3791] = "test_data_3791.txt";
test_data_files[3792] = "test_data_3792.txt";
test_data_files[3793] = "test_data_3793.txt";
test_data_files[3794] = "test_data_3794.txt";
test_data_files[3795] = "test_data_3795.txt";
test_data_files[3796] = "test_data_3796.txt";
test_data_files[3797] = "test_data_3797.txt";
test_data_files[3798] = "test_data_3798.txt";
test_data_files[3799] = "test_data_3799.txt";
test_data_files[3800] = "test_data_3800.txt";
test_data_files[3801] = "test_data_3801.txt";
test_data_files[3802] = "test_data_3802.txt";
test_data_files[3803] = "test_data_3803.txt";
test_data_files[3804] = "test_data_3804.txt";
test_data_files[3805] = "test_data_3805.txt";
test_data_files[3806] = "test_data_3806.txt";
test_data_files[3807] = "test_data_3807.txt";
test_data_files[3808] = "test_data_3808.txt";
test_data_files[3809] = "test_data_3809.txt";
test_data_files[3810] = "test_data_3810.txt";
test_data_files[3811] = "test_data_3811.txt";
test_data_files[3812] = "test_data_3812.txt";
test_data_files[3813] = "test_data_3813.txt";
test_data_files[3814] = "test_data_3814.txt";
test_data_files[3815] = "test_data_3815.txt";
test_data_files[3816] = "test_data_3816.txt";
test_data_files[3817] = "test_data_3817.txt";
test_data_files[3818] = "test_data_3818.txt";
test_data_files[3819] = "test_data_3819.txt";
test_data_files[3820] = "test_data_3820.txt";
test_data_files[3821] = "test_data_3821.txt";
test_data_files[3822] = "test_data_3822.txt";
test_data_files[3823] = "test_data_3823.txt";
test_data_files[3824] = "test_data_3824.txt";
test_data_files[3825] = "test_data_3825.txt";
test_data_files[3826] = "test_data_3826.txt";
test_data_files[3827] = "test_data_3827.txt";
test_data_files[3828] = "test_data_3828.txt";
test_data_files[3829] = "test_data_3829.txt";
test_data_files[3830] = "test_data_3830.txt";
test_data_files[3831] = "test_data_3831.txt";
test_data_files[3832] = "test_data_3832.txt";
test_data_files[3833] = "test_data_3833.txt";
test_data_files[3834] = "test_data_3834.txt";
test_data_files[3835] = "test_data_3835.txt";
test_data_files[3836] = "test_data_3836.txt";
test_data_files[3837] = "test_data_3837.txt";
test_data_files[3838] = "test_data_3838.txt";
test_data_files[3839] = "test_data_3839.txt";
test_data_files[3840] = "test_data_3840.txt";
test_data_files[3841] = "test_data_3841.txt";
test_data_files[3842] = "test_data_3842.txt";
test_data_files[3843] = "test_data_3843.txt";
test_data_files[3844] = "test_data_3844.txt";
test_data_files[3845] = "test_data_3845.txt";
test_data_files[3846] = "test_data_3846.txt";
test_data_files[3847] = "test_data_3847.txt";
test_data_files[3848] = "test_data_3848.txt";
test_data_files[3849] = "test_data_3849.txt";
test_data_files[3850] = "test_data_3850.txt";
test_data_files[3851] = "test_data_3851.txt";
test_data_files[3852] = "test_data_3852.txt";
test_data_files[3853] = "test_data_3853.txt";
test_data_files[3854] = "test_data_3854.txt";
test_data_files[3855] = "test_data_3855.txt";
test_data_files[3856] = "test_data_3856.txt";
test_data_files[3857] = "test_data_3857.txt";
test_data_files[3858] = "test_data_3858.txt";
test_data_files[3859] = "test_data_3859.txt";
test_data_files[3860] = "test_data_3860.txt";
test_data_files[3861] = "test_data_3861.txt";
test_data_files[3862] = "test_data_3862.txt";
test_data_files[3863] = "test_data_3863.txt";
test_data_files[3864] = "test_data_3864.txt";
test_data_files[3865] = "test_data_3865.txt";
test_data_files[3866] = "test_data_3866.txt";
test_data_files[3867] = "test_data_3867.txt";
test_data_files[3868] = "test_data_3868.txt";
test_data_files[3869] = "test_data_3869.txt";
test_data_files[3870] = "test_data_3870.txt";
test_data_files[3871] = "test_data_3871.txt";
test_data_files[3872] = "test_data_3872.txt";
test_data_files[3873] = "test_data_3873.txt";
test_data_files[3874] = "test_data_3874.txt";
test_data_files[3875] = "test_data_3875.txt";
test_data_files[3876] = "test_data_3876.txt";
test_data_files[3877] = "test_data_3877.txt";
test_data_files[3878] = "test_data_3878.txt";
test_data_files[3879] = "test_data_3879.txt";
test_data_files[3880] = "test_data_3880.txt";
test_data_files[3881] = "test_data_3881.txt";
test_data_files[3882] = "test_data_3882.txt";
test_data_files[3883] = "test_data_3883.txt";
test_data_files[3884] = "test_data_3884.txt";
test_data_files[3885] = "test_data_3885.txt";
test_data_files[3886] = "test_data_3886.txt";
test_data_files[3887] = "test_data_3887.txt";
test_data_files[3888] = "test_data_3888.txt";
test_data_files[3889] = "test_data_3889.txt";
test_data_files[3890] = "test_data_3890.txt";
test_data_files[3891] = "test_data_3891.txt";
test_data_files[3892] = "test_data_3892.txt";
test_data_files[3893] = "test_data_3893.txt";
test_data_files[3894] = "test_data_3894.txt";
test_data_files[3895] = "test_data_3895.txt";
test_data_files[3896] = "test_data_3896.txt";
test_data_files[3897] = "test_data_3897.txt";
test_data_files[3898] = "test_data_3898.txt";
test_data_files[3899] = "test_data_3899.txt";
test_data_files[3900] = "test_data_3900.txt";
test_data_files[3901] = "test_data_3901.txt";
test_data_files[3902] = "test_data_3902.txt";
test_data_files[3903] = "test_data_3903.txt";
test_data_files[3904] = "test_data_3904.txt";
test_data_files[3905] = "test_data_3905.txt";
test_data_files[3906] = "test_data_3906.txt";
test_data_files[3907] = "test_data_3907.txt";
test_data_files[3908] = "test_data_3908.txt";
test_data_files[3909] = "test_data_3909.txt";
test_data_files[3910] = "test_data_3910.txt";
test_data_files[3911] = "test_data_3911.txt";
test_data_files[3912] = "test_data_3912.txt";
test_data_files[3913] = "test_data_3913.txt";
test_data_files[3914] = "test_data_3914.txt";
test_data_files[3915] = "test_data_3915.txt";
test_data_files[3916] = "test_data_3916.txt";
test_data_files[3917] = "test_data_3917.txt";
test_data_files[3918] = "test_data_3918.txt";
test_data_files[3919] = "test_data_3919.txt";
test_data_files[3920] = "test_data_3920.txt";
test_data_files[3921] = "test_data_3921.txt";
test_data_files[3922] = "test_data_3922.txt";
test_data_files[3923] = "test_data_3923.txt";
test_data_files[3924] = "test_data_3924.txt";
test_data_files[3925] = "test_data_3925.txt";
test_data_files[3926] = "test_data_3926.txt";
test_data_files[3927] = "test_data_3927.txt";
test_data_files[3928] = "test_data_3928.txt";
test_data_files[3929] = "test_data_3929.txt";
test_data_files[3930] = "test_data_3930.txt";
test_data_files[3931] = "test_data_3931.txt";
test_data_files[3932] = "test_data_3932.txt";
test_data_files[3933] = "test_data_3933.txt";
test_data_files[3934] = "test_data_3934.txt";
test_data_files[3935] = "test_data_3935.txt";
test_data_files[3936] = "test_data_3936.txt";
test_data_files[3937] = "test_data_3937.txt";
test_data_files[3938] = "test_data_3938.txt";
test_data_files[3939] = "test_data_3939.txt";
test_data_files[3940] = "test_data_3940.txt";
test_data_files[3941] = "test_data_3941.txt";
test_data_files[3942] = "test_data_3942.txt";
test_data_files[3943] = "test_data_3943.txt";
test_data_files[3944] = "test_data_3944.txt";
test_data_files[3945] = "test_data_3945.txt";
test_data_files[3946] = "test_data_3946.txt";
test_data_files[3947] = "test_data_3947.txt";
test_data_files[3948] = "test_data_3948.txt";
test_data_files[3949] = "test_data_3949.txt";
test_data_files[3950] = "test_data_3950.txt";
test_data_files[3951] = "test_data_3951.txt";
test_data_files[3952] = "test_data_3952.txt";
test_data_files[3953] = "test_data_3953.txt";
test_data_files[3954] = "test_data_3954.txt";
test_data_files[3955] = "test_data_3955.txt";
test_data_files[3956] = "test_data_3956.txt";
test_data_files[3957] = "test_data_3957.txt";
test_data_files[3958] = "test_data_3958.txt";
test_data_files[3959] = "test_data_3959.txt";
test_data_files[3960] = "test_data_3960.txt";
test_data_files[3961] = "test_data_3961.txt";
test_data_files[3962] = "test_data_3962.txt";
test_data_files[3963] = "test_data_3963.txt";
test_data_files[3964] = "test_data_3964.txt";
test_data_files[3965] = "test_data_3965.txt";
test_data_files[3966] = "test_data_3966.txt";
test_data_files[3967] = "test_data_3967.txt";
test_data_files[3968] = "test_data_3968.txt";
test_data_files[3969] = "test_data_3969.txt";
test_data_files[3970] = "test_data_3970.txt";
test_data_files[3971] = "test_data_3971.txt";
test_data_files[3972] = "test_data_3972.txt";
test_data_files[3973] = "test_data_3973.txt";
test_data_files[3974] = "test_data_3974.txt";
test_data_files[3975] = "test_data_3975.txt";
test_data_files[3976] = "test_data_3976.txt";
test_data_files[3977] = "test_data_3977.txt";
test_data_files[3978] = "test_data_3978.txt";
test_data_files[3979] = "test_data_3979.txt";
test_data_files[3980] = "test_data_3980.txt";
test_data_files[3981] = "test_data_3981.txt";
test_data_files[3982] = "test_data_3982.txt";
test_data_files[3983] = "test_data_3983.txt";
test_data_files[3984] = "test_data_3984.txt";
test_data_files[3985] = "test_data_3985.txt";
test_data_files[3986] = "test_data_3986.txt";
test_data_files[3987] = "test_data_3987.txt";
test_data_files[3988] = "test_data_3988.txt";
test_data_files[3989] = "test_data_3989.txt";
test_data_files[3990] = "test_data_3990.txt";
test_data_files[3991] = "test_data_3991.txt";
test_data_files[3992] = "test_data_3992.txt";
test_data_files[3993] = "test_data_3993.txt";
test_data_files[3994] = "test_data_3994.txt";
test_data_files[3995] = "test_data_3995.txt";
test_data_files[3996] = "test_data_3996.txt";
test_data_files[3997] = "test_data_3997.txt";
test_data_files[3998] = "test_data_3998.txt";
test_data_files[3999] = "test_data_3999.txt";
test_data_files[4000] = "test_data_4000.txt";
test_data_files[4001] = "test_data_4001.txt";
test_data_files[4002] = "test_data_4002.txt";
test_data_files[4003] = "test_data_4003.txt";
test_data_files[4004] = "test_data_4004.txt";
test_data_files[4005] = "test_data_4005.txt";
test_data_files[4006] = "test_data_4006.txt";
test_data_files[4007] = "test_data_4007.txt";
test_data_files[4008] = "test_data_4008.txt";
test_data_files[4009] = "test_data_4009.txt";
test_data_files[4010] = "test_data_4010.txt";
test_data_files[4011] = "test_data_4011.txt";
test_data_files[4012] = "test_data_4012.txt";
test_data_files[4013] = "test_data_4013.txt";
test_data_files[4014] = "test_data_4014.txt";
test_data_files[4015] = "test_data_4015.txt";
test_data_files[4016] = "test_data_4016.txt";
test_data_files[4017] = "test_data_4017.txt";
test_data_files[4018] = "test_data_4018.txt";
test_data_files[4019] = "test_data_4019.txt";
test_data_files[4020] = "test_data_4020.txt";
test_data_files[4021] = "test_data_4021.txt";
test_data_files[4022] = "test_data_4022.txt";
test_data_files[4023] = "test_data_4023.txt";
test_data_files[4024] = "test_data_4024.txt";
test_data_files[4025] = "test_data_4025.txt";
test_data_files[4026] = "test_data_4026.txt";
test_data_files[4027] = "test_data_4027.txt";
test_data_files[4028] = "test_data_4028.txt";
test_data_files[4029] = "test_data_4029.txt";
test_data_files[4030] = "test_data_4030.txt";
test_data_files[4031] = "test_data_4031.txt";
test_data_files[4032] = "test_data_4032.txt";
test_data_files[4033] = "test_data_4033.txt";
test_data_files[4034] = "test_data_4034.txt";
test_data_files[4035] = "test_data_4035.txt";
test_data_files[4036] = "test_data_4036.txt";
test_data_files[4037] = "test_data_4037.txt";
test_data_files[4038] = "test_data_4038.txt";
test_data_files[4039] = "test_data_4039.txt";
test_data_files[4040] = "test_data_4040.txt";
test_data_files[4041] = "test_data_4041.txt";
test_data_files[4042] = "test_data_4042.txt";
test_data_files[4043] = "test_data_4043.txt";
test_data_files[4044] = "test_data_4044.txt";
test_data_files[4045] = "test_data_4045.txt";
test_data_files[4046] = "test_data_4046.txt";
test_data_files[4047] = "test_data_4047.txt";
test_data_files[4048] = "test_data_4048.txt";
test_data_files[4049] = "test_data_4049.txt";
test_data_files[4050] = "test_data_4050.txt";
test_data_files[4051] = "test_data_4051.txt";
test_data_files[4052] = "test_data_4052.txt";
test_data_files[4053] = "test_data_4053.txt";
test_data_files[4054] = "test_data_4054.txt";
test_data_files[4055] = "test_data_4055.txt";
test_data_files[4056] = "test_data_4056.txt";
test_data_files[4057] = "test_data_4057.txt";
test_data_files[4058] = "test_data_4058.txt";
test_data_files[4059] = "test_data_4059.txt";
test_data_files[4060] = "test_data_4060.txt";
test_data_files[4061] = "test_data_4061.txt";
test_data_files[4062] = "test_data_4062.txt";
test_data_files[4063] = "test_data_4063.txt";
test_data_files[4064] = "test_data_4064.txt";
test_data_files[4065] = "test_data_4065.txt";
test_data_files[4066] = "test_data_4066.txt";
test_data_files[4067] = "test_data_4067.txt";
test_data_files[4068] = "test_data_4068.txt";
test_data_files[4069] = "test_data_4069.txt";
test_data_files[4070] = "test_data_4070.txt";
test_data_files[4071] = "test_data_4071.txt";
test_data_files[4072] = "test_data_4072.txt";
test_data_files[4073] = "test_data_4073.txt";
test_data_files[4074] = "test_data_4074.txt";
test_data_files[4075] = "test_data_4075.txt";
test_data_files[4076] = "test_data_4076.txt";
test_data_files[4077] = "test_data_4077.txt";
test_data_files[4078] = "test_data_4078.txt";
test_data_files[4079] = "test_data_4079.txt";
test_data_files[4080] = "test_data_4080.txt";
test_data_files[4081] = "test_data_4081.txt";
test_data_files[4082] = "test_data_4082.txt";
test_data_files[4083] = "test_data_4083.txt";
test_data_files[4084] = "test_data_4084.txt";
test_data_files[4085] = "test_data_4085.txt";
test_data_files[4086] = "test_data_4086.txt";
test_data_files[4087] = "test_data_4087.txt";
test_data_files[4088] = "test_data_4088.txt";
test_data_files[4089] = "test_data_4089.txt";
test_data_files[4090] = "test_data_4090.txt";
test_data_files[4091] = "test_data_4091.txt";
test_data_files[4092] = "test_data_4092.txt";
test_data_files[4093] = "test_data_4093.txt";
test_data_files[4094] = "test_data_4094.txt";
test_data_files[4095] = "test_data_4095.txt";
test_data_files[4096] = "test_data_4096.txt";
test_data_files[4097] = "test_data_4097.txt";
test_data_files[4098] = "test_data_4098.txt";
test_data_files[4099] = "test_data_4099.txt";
test_data_files[4100] = "test_data_4100.txt";
test_data_files[4101] = "test_data_4101.txt";
test_data_files[4102] = "test_data_4102.txt";
test_data_files[4103] = "test_data_4103.txt";
test_data_files[4104] = "test_data_4104.txt";
test_data_files[4105] = "test_data_4105.txt";
test_data_files[4106] = "test_data_4106.txt";
test_data_files[4107] = "test_data_4107.txt";
test_data_files[4108] = "test_data_4108.txt";
test_data_files[4109] = "test_data_4109.txt";
test_data_files[4110] = "test_data_4110.txt";
test_data_files[4111] = "test_data_4111.txt";
test_data_files[4112] = "test_data_4112.txt";
test_data_files[4113] = "test_data_4113.txt";
test_data_files[4114] = "test_data_4114.txt";
test_data_files[4115] = "test_data_4115.txt";
test_data_files[4116] = "test_data_4116.txt";
test_data_files[4117] = "test_data_4117.txt";
test_data_files[4118] = "test_data_4118.txt";
test_data_files[4119] = "test_data_4119.txt";
test_data_files[4120] = "test_data_4120.txt";
test_data_files[4121] = "test_data_4121.txt";
test_data_files[4122] = "test_data_4122.txt";
test_data_files[4123] = "test_data_4123.txt";
test_data_files[4124] = "test_data_4124.txt";
test_data_files[4125] = "test_data_4125.txt";
test_data_files[4126] = "test_data_4126.txt";
test_data_files[4127] = "test_data_4127.txt";
test_data_files[4128] = "test_data_4128.txt";
test_data_files[4129] = "test_data_4129.txt";
test_data_files[4130] = "test_data_4130.txt";
test_data_files[4131] = "test_data_4131.txt";
test_data_files[4132] = "test_data_4132.txt";
test_data_files[4133] = "test_data_4133.txt";
test_data_files[4134] = "test_data_4134.txt";
test_data_files[4135] = "test_data_4135.txt";
test_data_files[4136] = "test_data_4136.txt";
test_data_files[4137] = "test_data_4137.txt";
test_data_files[4138] = "test_data_4138.txt";
test_data_files[4139] = "test_data_4139.txt";
test_data_files[4140] = "test_data_4140.txt";
test_data_files[4141] = "test_data_4141.txt";
test_data_files[4142] = "test_data_4142.txt";
test_data_files[4143] = "test_data_4143.txt";
test_data_files[4144] = "test_data_4144.txt";
test_data_files[4145] = "test_data_4145.txt";
test_data_files[4146] = "test_data_4146.txt";
test_data_files[4147] = "test_data_4147.txt";
test_data_files[4148] = "test_data_4148.txt";
test_data_files[4149] = "test_data_4149.txt";
test_data_files[4150] = "test_data_4150.txt";
test_data_files[4151] = "test_data_4151.txt";
test_data_files[4152] = "test_data_4152.txt";
test_data_files[4153] = "test_data_4153.txt";
test_data_files[4154] = "test_data_4154.txt";
test_data_files[4155] = "test_data_4155.txt";
test_data_files[4156] = "test_data_4156.txt";
test_data_files[4157] = "test_data_4157.txt";
test_data_files[4158] = "test_data_4158.txt";
test_data_files[4159] = "test_data_4159.txt";
test_data_files[4160] = "test_data_4160.txt";
test_data_files[4161] = "test_data_4161.txt";
test_data_files[4162] = "test_data_4162.txt";
test_data_files[4163] = "test_data_4163.txt";
test_data_files[4164] = "test_data_4164.txt";
test_data_files[4165] = "test_data_4165.txt";
test_data_files[4166] = "test_data_4166.txt";
test_data_files[4167] = "test_data_4167.txt";
test_data_files[4168] = "test_data_4168.txt";
test_data_files[4169] = "test_data_4169.txt";
test_data_files[4170] = "test_data_4170.txt";
test_data_files[4171] = "test_data_4171.txt";
test_data_files[4172] = "test_data_4172.txt";
test_data_files[4173] = "test_data_4173.txt";
test_data_files[4174] = "test_data_4174.txt";
test_data_files[4175] = "test_data_4175.txt";
test_data_files[4176] = "test_data_4176.txt";
test_data_files[4177] = "test_data_4177.txt";
test_data_files[4178] = "test_data_4178.txt";
test_data_files[4179] = "test_data_4179.txt";
test_data_files[4180] = "test_data_4180.txt";
test_data_files[4181] = "test_data_4181.txt";
test_data_files[4182] = "test_data_4182.txt";
test_data_files[4183] = "test_data_4183.txt";
test_data_files[4184] = "test_data_4184.txt";
test_data_files[4185] = "test_data_4185.txt";
test_data_files[4186] = "test_data_4186.txt";
test_data_files[4187] = "test_data_4187.txt";
test_data_files[4188] = "test_data_4188.txt";
test_data_files[4189] = "test_data_4189.txt";
test_data_files[4190] = "test_data_4190.txt";
test_data_files[4191] = "test_data_4191.txt";
test_data_files[4192] = "test_data_4192.txt";
test_data_files[4193] = "test_data_4193.txt";
test_data_files[4194] = "test_data_4194.txt";
test_data_files[4195] = "test_data_4195.txt";
test_data_files[4196] = "test_data_4196.txt";
test_data_files[4197] = "test_data_4197.txt";
test_data_files[4198] = "test_data_4198.txt";
test_data_files[4199] = "test_data_4199.txt";
test_data_files[4200] = "test_data_4200.txt";
test_data_files[4201] = "test_data_4201.txt";
test_data_files[4202] = "test_data_4202.txt";
test_data_files[4203] = "test_data_4203.txt";
test_data_files[4204] = "test_data_4204.txt";
test_data_files[4205] = "test_data_4205.txt";
test_data_files[4206] = "test_data_4206.txt";
test_data_files[4207] = "test_data_4207.txt";
test_data_files[4208] = "test_data_4208.txt";
test_data_files[4209] = "test_data_4209.txt";
test_data_files[4210] = "test_data_4210.txt";
test_data_files[4211] = "test_data_4211.txt";
test_data_files[4212] = "test_data_4212.txt";
test_data_files[4213] = "test_data_4213.txt";
test_data_files[4214] = "test_data_4214.txt";
test_data_files[4215] = "test_data_4215.txt";
test_data_files[4216] = "test_data_4216.txt";
test_data_files[4217] = "test_data_4217.txt";
test_data_files[4218] = "test_data_4218.txt";
test_data_files[4219] = "test_data_4219.txt";
test_data_files[4220] = "test_data_4220.txt";
test_data_files[4221] = "test_data_4221.txt";
test_data_files[4222] = "test_data_4222.txt";
test_data_files[4223] = "test_data_4223.txt";
test_data_files[4224] = "test_data_4224.txt";
test_data_files[4225] = "test_data_4225.txt";
test_data_files[4226] = "test_data_4226.txt";
test_data_files[4227] = "test_data_4227.txt";
test_data_files[4228] = "test_data_4228.txt";
test_data_files[4229] = "test_data_4229.txt";
test_data_files[4230] = "test_data_4230.txt";
test_data_files[4231] = "test_data_4231.txt";
test_data_files[4232] = "test_data_4232.txt";
test_data_files[4233] = "test_data_4233.txt";
test_data_files[4234] = "test_data_4234.txt";
test_data_files[4235] = "test_data_4235.txt";
test_data_files[4236] = "test_data_4236.txt";
test_data_files[4237] = "test_data_4237.txt";
test_data_files[4238] = "test_data_4238.txt";
test_data_files[4239] = "test_data_4239.txt";
test_data_files[4240] = "test_data_4240.txt";
test_data_files[4241] = "test_data_4241.txt";
test_data_files[4242] = "test_data_4242.txt";
test_data_files[4243] = "test_data_4243.txt";
test_data_files[4244] = "test_data_4244.txt";
test_data_files[4245] = "test_data_4245.txt";
test_data_files[4246] = "test_data_4246.txt";
test_data_files[4247] = "test_data_4247.txt";
test_data_files[4248] = "test_data_4248.txt";
test_data_files[4249] = "test_data_4249.txt";
test_data_files[4250] = "test_data_4250.txt";
test_data_files[4251] = "test_data_4251.txt";
test_data_files[4252] = "test_data_4252.txt";
test_data_files[4253] = "test_data_4253.txt";
test_data_files[4254] = "test_data_4254.txt";
test_data_files[4255] = "test_data_4255.txt";
test_data_files[4256] = "test_data_4256.txt";
test_data_files[4257] = "test_data_4257.txt";
test_data_files[4258] = "test_data_4258.txt";
test_data_files[4259] = "test_data_4259.txt";
test_data_files[4260] = "test_data_4260.txt";
test_data_files[4261] = "test_data_4261.txt";
test_data_files[4262] = "test_data_4262.txt";
test_data_files[4263] = "test_data_4263.txt";
test_data_files[4264] = "test_data_4264.txt";
test_data_files[4265] = "test_data_4265.txt";
test_data_files[4266] = "test_data_4266.txt";
test_data_files[4267] = "test_data_4267.txt";
test_data_files[4268] = "test_data_4268.txt";
test_data_files[4269] = "test_data_4269.txt";
test_data_files[4270] = "test_data_4270.txt";
test_data_files[4271] = "test_data_4271.txt";
test_data_files[4272] = "test_data_4272.txt";
test_data_files[4273] = "test_data_4273.txt";
test_data_files[4274] = "test_data_4274.txt";
test_data_files[4275] = "test_data_4275.txt";
test_data_files[4276] = "test_data_4276.txt";
test_data_files[4277] = "test_data_4277.txt";
test_data_files[4278] = "test_data_4278.txt";
test_data_files[4279] = "test_data_4279.txt";
test_data_files[4280] = "test_data_4280.txt";
test_data_files[4281] = "test_data_4281.txt";
test_data_files[4282] = "test_data_4282.txt";
test_data_files[4283] = "test_data_4283.txt";
test_data_files[4284] = "test_data_4284.txt";
test_data_files[4285] = "test_data_4285.txt";
test_data_files[4286] = "test_data_4286.txt";
test_data_files[4287] = "test_data_4287.txt";
test_data_files[4288] = "test_data_4288.txt";
test_data_files[4289] = "test_data_4289.txt";
test_data_files[4290] = "test_data_4290.txt";
test_data_files[4291] = "test_data_4291.txt";
test_data_files[4292] = "test_data_4292.txt";
test_data_files[4293] = "test_data_4293.txt";
test_data_files[4294] = "test_data_4294.txt";
test_data_files[4295] = "test_data_4295.txt";
test_data_files[4296] = "test_data_4296.txt";
test_data_files[4297] = "test_data_4297.txt";
test_data_files[4298] = "test_data_4298.txt";
test_data_files[4299] = "test_data_4299.txt";
test_data_files[4300] = "test_data_4300.txt";
test_data_files[4301] = "test_data_4301.txt";
test_data_files[4302] = "test_data_4302.txt";
test_data_files[4303] = "test_data_4303.txt";
test_data_files[4304] = "test_data_4304.txt";
test_data_files[4305] = "test_data_4305.txt";
test_data_files[4306] = "test_data_4306.txt";
test_data_files[4307] = "test_data_4307.txt";
test_data_files[4308] = "test_data_4308.txt";
test_data_files[4309] = "test_data_4309.txt";
test_data_files[4310] = "test_data_4310.txt";
test_data_files[4311] = "test_data_4311.txt";
test_data_files[4312] = "test_data_4312.txt";
test_data_files[4313] = "test_data_4313.txt";
test_data_files[4314] = "test_data_4314.txt";
test_data_files[4315] = "test_data_4315.txt";
test_data_files[4316] = "test_data_4316.txt";
test_data_files[4317] = "test_data_4317.txt";
test_data_files[4318] = "test_data_4318.txt";
test_data_files[4319] = "test_data_4319.txt";
test_data_files[4320] = "test_data_4320.txt";
test_data_files[4321] = "test_data_4321.txt";
test_data_files[4322] = "test_data_4322.txt";
test_data_files[4323] = "test_data_4323.txt";
test_data_files[4324] = "test_data_4324.txt";
test_data_files[4325] = "test_data_4325.txt";
test_data_files[4326] = "test_data_4326.txt";
test_data_files[4327] = "test_data_4327.txt";
test_data_files[4328] = "test_data_4328.txt";
test_data_files[4329] = "test_data_4329.txt";
test_data_files[4330] = "test_data_4330.txt";
test_data_files[4331] = "test_data_4331.txt";
test_data_files[4332] = "test_data_4332.txt";
test_data_files[4333] = "test_data_4333.txt";
test_data_files[4334] = "test_data_4334.txt";
test_data_files[4335] = "test_data_4335.txt";
test_data_files[4336] = "test_data_4336.txt";
test_data_files[4337] = "test_data_4337.txt";
test_data_files[4338] = "test_data_4338.txt";
test_data_files[4339] = "test_data_4339.txt";
test_data_files[4340] = "test_data_4340.txt";
test_data_files[4341] = "test_data_4341.txt";
test_data_files[4342] = "test_data_4342.txt";
test_data_files[4343] = "test_data_4343.txt";
test_data_files[4344] = "test_data_4344.txt";
test_data_files[4345] = "test_data_4345.txt";
test_data_files[4346] = "test_data_4346.txt";
test_data_files[4347] = "test_data_4347.txt";
test_data_files[4348] = "test_data_4348.txt";
test_data_files[4349] = "test_data_4349.txt";
test_data_files[4350] = "test_data_4350.txt";
test_data_files[4351] = "test_data_4351.txt";
test_data_files[4352] = "test_data_4352.txt";
test_data_files[4353] = "test_data_4353.txt";
test_data_files[4354] = "test_data_4354.txt";
test_data_files[4355] = "test_data_4355.txt";
test_data_files[4356] = "test_data_4356.txt";
test_data_files[4357] = "test_data_4357.txt";
test_data_files[4358] = "test_data_4358.txt";
test_data_files[4359] = "test_data_4359.txt";
test_data_files[4360] = "test_data_4360.txt";
test_data_files[4361] = "test_data_4361.txt";
test_data_files[4362] = "test_data_4362.txt";
test_data_files[4363] = "test_data_4363.txt";
test_data_files[4364] = "test_data_4364.txt";
test_data_files[4365] = "test_data_4365.txt";
test_data_files[4366] = "test_data_4366.txt";
test_data_files[4367] = "test_data_4367.txt";
test_data_files[4368] = "test_data_4368.txt";
test_data_files[4369] = "test_data_4369.txt";
test_data_files[4370] = "test_data_4370.txt";
test_data_files[4371] = "test_data_4371.txt";
test_data_files[4372] = "test_data_4372.txt";
test_data_files[4373] = "test_data_4373.txt";
test_data_files[4374] = "test_data_4374.txt";
test_data_files[4375] = "test_data_4375.txt";
test_data_files[4376] = "test_data_4376.txt";
test_data_files[4377] = "test_data_4377.txt";
test_data_files[4378] = "test_data_4378.txt";
test_data_files[4379] = "test_data_4379.txt";
test_data_files[4380] = "test_data_4380.txt";
test_data_files[4381] = "test_data_4381.txt";
test_data_files[4382] = "test_data_4382.txt";
test_data_files[4383] = "test_data_4383.txt";
test_data_files[4384] = "test_data_4384.txt";
test_data_files[4385] = "test_data_4385.txt";
test_data_files[4386] = "test_data_4386.txt";
test_data_files[4387] = "test_data_4387.txt";
test_data_files[4388] = "test_data_4388.txt";
test_data_files[4389] = "test_data_4389.txt";
test_data_files[4390] = "test_data_4390.txt";
test_data_files[4391] = "test_data_4391.txt";
test_data_files[4392] = "test_data_4392.txt";
test_data_files[4393] = "test_data_4393.txt";
test_data_files[4394] = "test_data_4394.txt";
test_data_files[4395] = "test_data_4395.txt";
test_data_files[4396] = "test_data_4396.txt";
test_data_files[4397] = "test_data_4397.txt";
test_data_files[4398] = "test_data_4398.txt";
test_data_files[4399] = "test_data_4399.txt";
test_data_files[4400] = "test_data_4400.txt";
test_data_files[4401] = "test_data_4401.txt";
test_data_files[4402] = "test_data_4402.txt";
test_data_files[4403] = "test_data_4403.txt";
test_data_files[4404] = "test_data_4404.txt";
test_data_files[4405] = "test_data_4405.txt";
test_data_files[4406] = "test_data_4406.txt";
test_data_files[4407] = "test_data_4407.txt";
test_data_files[4408] = "test_data_4408.txt";
test_data_files[4409] = "test_data_4409.txt";
test_data_files[4410] = "test_data_4410.txt";
test_data_files[4411] = "test_data_4411.txt";
test_data_files[4412] = "test_data_4412.txt";
test_data_files[4413] = "test_data_4413.txt";
test_data_files[4414] = "test_data_4414.txt";
test_data_files[4415] = "test_data_4415.txt";
test_data_files[4416] = "test_data_4416.txt";
test_data_files[4417] = "test_data_4417.txt";
test_data_files[4418] = "test_data_4418.txt";
test_data_files[4419] = "test_data_4419.txt";
test_data_files[4420] = "test_data_4420.txt";
test_data_files[4421] = "test_data_4421.txt";
test_data_files[4422] = "test_data_4422.txt";
test_data_files[4423] = "test_data_4423.txt";
test_data_files[4424] = "test_data_4424.txt";
test_data_files[4425] = "test_data_4425.txt";
test_data_files[4426] = "test_data_4426.txt";
test_data_files[4427] = "test_data_4427.txt";
test_data_files[4428] = "test_data_4428.txt";
test_data_files[4429] = "test_data_4429.txt";
test_data_files[4430] = "test_data_4430.txt";
test_data_files[4431] = "test_data_4431.txt";
test_data_files[4432] = "test_data_4432.txt";
test_data_files[4433] = "test_data_4433.txt";
test_data_files[4434] = "test_data_4434.txt";
test_data_files[4435] = "test_data_4435.txt";
test_data_files[4436] = "test_data_4436.txt";
test_data_files[4437] = "test_data_4437.txt";
test_data_files[4438] = "test_data_4438.txt";
test_data_files[4439] = "test_data_4439.txt";
test_data_files[4440] = "test_data_4440.txt";
test_data_files[4441] = "test_data_4441.txt";
test_data_files[4442] = "test_data_4442.txt";
test_data_files[4443] = "test_data_4443.txt";
test_data_files[4444] = "test_data_4444.txt";
test_data_files[4445] = "test_data_4445.txt";
test_data_files[4446] = "test_data_4446.txt";
test_data_files[4447] = "test_data_4447.txt";
test_data_files[4448] = "test_data_4448.txt";
test_data_files[4449] = "test_data_4449.txt";
test_data_files[4450] = "test_data_4450.txt";
test_data_files[4451] = "test_data_4451.txt";
test_data_files[4452] = "test_data_4452.txt";
test_data_files[4453] = "test_data_4453.txt";
test_data_files[4454] = "test_data_4454.txt";
test_data_files[4455] = "test_data_4455.txt";
test_data_files[4456] = "test_data_4456.txt";
test_data_files[4457] = "test_data_4457.txt";
test_data_files[4458] = "test_data_4458.txt";
test_data_files[4459] = "test_data_4459.txt";
test_data_files[4460] = "test_data_4460.txt";
test_data_files[4461] = "test_data_4461.txt";
test_data_files[4462] = "test_data_4462.txt";
test_data_files[4463] = "test_data_4463.txt";
test_data_files[4464] = "test_data_4464.txt";
test_data_files[4465] = "test_data_4465.txt";
test_data_files[4466] = "test_data_4466.txt";
test_data_files[4467] = "test_data_4467.txt";
test_data_files[4468] = "test_data_4468.txt";
test_data_files[4469] = "test_data_4469.txt";
test_data_files[4470] = "test_data_4470.txt";
test_data_files[4471] = "test_data_4471.txt";
test_data_files[4472] = "test_data_4472.txt";
test_data_files[4473] = "test_data_4473.txt";
test_data_files[4474] = "test_data_4474.txt";
test_data_files[4475] = "test_data_4475.txt";
test_data_files[4476] = "test_data_4476.txt";
test_data_files[4477] = "test_data_4477.txt";
test_data_files[4478] = "test_data_4478.txt";
test_data_files[4479] = "test_data_4479.txt";
test_data_files[4480] = "test_data_4480.txt";
test_data_files[4481] = "test_data_4481.txt";
test_data_files[4482] = "test_data_4482.txt";
test_data_files[4483] = "test_data_4483.txt";
test_data_files[4484] = "test_data_4484.txt";
test_data_files[4485] = "test_data_4485.txt";
test_data_files[4486] = "test_data_4486.txt";
test_data_files[4487] = "test_data_4487.txt";
test_data_files[4488] = "test_data_4488.txt";
test_data_files[4489] = "test_data_4489.txt";
test_data_files[4490] = "test_data_4490.txt";
test_data_files[4491] = "test_data_4491.txt";
test_data_files[4492] = "test_data_4492.txt";
test_data_files[4493] = "test_data_4493.txt";
test_data_files[4494] = "test_data_4494.txt";
test_data_files[4495] = "test_data_4495.txt";
test_data_files[4496] = "test_data_4496.txt";
test_data_files[4497] = "test_data_4497.txt";
test_data_files[4498] = "test_data_4498.txt";
test_data_files[4499] = "test_data_4499.txt";
test_data_files[4500] = "test_data_4500.txt";
test_data_files[4501] = "test_data_4501.txt";
test_data_files[4502] = "test_data_4502.txt";
test_data_files[4503] = "test_data_4503.txt";
test_data_files[4504] = "test_data_4504.txt";
test_data_files[4505] = "test_data_4505.txt";
test_data_files[4506] = "test_data_4506.txt";
test_data_files[4507] = "test_data_4507.txt";
test_data_files[4508] = "test_data_4508.txt";
test_data_files[4509] = "test_data_4509.txt";
test_data_files[4510] = "test_data_4510.txt";
test_data_files[4511] = "test_data_4511.txt";
test_data_files[4512] = "test_data_4512.txt";
test_data_files[4513] = "test_data_4513.txt";
test_data_files[4514] = "test_data_4514.txt";
test_data_files[4515] = "test_data_4515.txt";
test_data_files[4516] = "test_data_4516.txt";
test_data_files[4517] = "test_data_4517.txt";
test_data_files[4518] = "test_data_4518.txt";
test_data_files[4519] = "test_data_4519.txt";
test_data_files[4520] = "test_data_4520.txt";
test_data_files[4521] = "test_data_4521.txt";
test_data_files[4522] = "test_data_4522.txt";
test_data_files[4523] = "test_data_4523.txt";
test_data_files[4524] = "test_data_4524.txt";
test_data_files[4525] = "test_data_4525.txt";
test_data_files[4526] = "test_data_4526.txt";
test_data_files[4527] = "test_data_4527.txt";
test_data_files[4528] = "test_data_4528.txt";
test_data_files[4529] = "test_data_4529.txt";
test_data_files[4530] = "test_data_4530.txt";
test_data_files[4531] = "test_data_4531.txt";
test_data_files[4532] = "test_data_4532.txt";
test_data_files[4533] = "test_data_4533.txt";
test_data_files[4534] = "test_data_4534.txt";
test_data_files[4535] = "test_data_4535.txt";
test_data_files[4536] = "test_data_4536.txt";
test_data_files[4537] = "test_data_4537.txt";
test_data_files[4538] = "test_data_4538.txt";
test_data_files[4539] = "test_data_4539.txt";
test_data_files[4540] = "test_data_4540.txt";
test_data_files[4541] = "test_data_4541.txt";
test_data_files[4542] = "test_data_4542.txt";
test_data_files[4543] = "test_data_4543.txt";
test_data_files[4544] = "test_data_4544.txt";
test_data_files[4545] = "test_data_4545.txt";
test_data_files[4546] = "test_data_4546.txt";
test_data_files[4547] = "test_data_4547.txt";
test_data_files[4548] = "test_data_4548.txt";
test_data_files[4549] = "test_data_4549.txt";
test_data_files[4550] = "test_data_4550.txt";
test_data_files[4551] = "test_data_4551.txt";
test_data_files[4552] = "test_data_4552.txt";
test_data_files[4553] = "test_data_4553.txt";
test_data_files[4554] = "test_data_4554.txt";
test_data_files[4555] = "test_data_4555.txt";
test_data_files[4556] = "test_data_4556.txt";
test_data_files[4557] = "test_data_4557.txt";
test_data_files[4558] = "test_data_4558.txt";
test_data_files[4559] = "test_data_4559.txt";
test_data_files[4560] = "test_data_4560.txt";
test_data_files[4561] = "test_data_4561.txt";
test_data_files[4562] = "test_data_4562.txt";
test_data_files[4563] = "test_data_4563.txt";
test_data_files[4564] = "test_data_4564.txt";
test_data_files[4565] = "test_data_4565.txt";
test_data_files[4566] = "test_data_4566.txt";
test_data_files[4567] = "test_data_4567.txt";
test_data_files[4568] = "test_data_4568.txt";
test_data_files[4569] = "test_data_4569.txt";
test_data_files[4570] = "test_data_4570.txt";
test_data_files[4571] = "test_data_4571.txt";
test_data_files[4572] = "test_data_4572.txt";
test_data_files[4573] = "test_data_4573.txt";
test_data_files[4574] = "test_data_4574.txt";
test_data_files[4575] = "test_data_4575.txt";
test_data_files[4576] = "test_data_4576.txt";
test_data_files[4577] = "test_data_4577.txt";
test_data_files[4578] = "test_data_4578.txt";
test_data_files[4579] = "test_data_4579.txt";
test_data_files[4580] = "test_data_4580.txt";
test_data_files[4581] = "test_data_4581.txt";
test_data_files[4582] = "test_data_4582.txt";
test_data_files[4583] = "test_data_4583.txt";
test_data_files[4584] = "test_data_4584.txt";
test_data_files[4585] = "test_data_4585.txt";
test_data_files[4586] = "test_data_4586.txt";
test_data_files[4587] = "test_data_4587.txt";
test_data_files[4588] = "test_data_4588.txt";
test_data_files[4589] = "test_data_4589.txt";
test_data_files[4590] = "test_data_4590.txt";
test_data_files[4591] = "test_data_4591.txt";
test_data_files[4592] = "test_data_4592.txt";
test_data_files[4593] = "test_data_4593.txt";
test_data_files[4594] = "test_data_4594.txt";
test_data_files[4595] = "test_data_4595.txt";
test_data_files[4596] = "test_data_4596.txt";
test_data_files[4597] = "test_data_4597.txt";
test_data_files[4598] = "test_data_4598.txt";
test_data_files[4599] = "test_data_4599.txt";
test_data_files[4600] = "test_data_4600.txt";
test_data_files[4601] = "test_data_4601.txt";
test_data_files[4602] = "test_data_4602.txt";
test_data_files[4603] = "test_data_4603.txt";
test_data_files[4604] = "test_data_4604.txt";
test_data_files[4605] = "test_data_4605.txt";
test_data_files[4606] = "test_data_4606.txt";
test_data_files[4607] = "test_data_4607.txt";
test_data_files[4608] = "test_data_4608.txt";
test_data_files[4609] = "test_data_4609.txt";
test_data_files[4610] = "test_data_4610.txt";
test_data_files[4611] = "test_data_4611.txt";
test_data_files[4612] = "test_data_4612.txt";
test_data_files[4613] = "test_data_4613.txt";
test_data_files[4614] = "test_data_4614.txt";
test_data_files[4615] = "test_data_4615.txt";
test_data_files[4616] = "test_data_4616.txt";
test_data_files[4617] = "test_data_4617.txt";
test_data_files[4618] = "test_data_4618.txt";
test_data_files[4619] = "test_data_4619.txt";
test_data_files[4620] = "test_data_4620.txt";
test_data_files[4621] = "test_data_4621.txt";
test_data_files[4622] = "test_data_4622.txt";
test_data_files[4623] = "test_data_4623.txt";
test_data_files[4624] = "test_data_4624.txt";
test_data_files[4625] = "test_data_4625.txt";
test_data_files[4626] = "test_data_4626.txt";
test_data_files[4627] = "test_data_4627.txt";
test_data_files[4628] = "test_data_4628.txt";
test_data_files[4629] = "test_data_4629.txt";
test_data_files[4630] = "test_data_4630.txt";
test_data_files[4631] = "test_data_4631.txt";
test_data_files[4632] = "test_data_4632.txt";
test_data_files[4633] = "test_data_4633.txt";
test_data_files[4634] = "test_data_4634.txt";
test_data_files[4635] = "test_data_4635.txt";
test_data_files[4636] = "test_data_4636.txt";
test_data_files[4637] = "test_data_4637.txt";
test_data_files[4638] = "test_data_4638.txt";
test_data_files[4639] = "test_data_4639.txt";
test_data_files[4640] = "test_data_4640.txt";
test_data_files[4641] = "test_data_4641.txt";
test_data_files[4642] = "test_data_4642.txt";
test_data_files[4643] = "test_data_4643.txt";
test_data_files[4644] = "test_data_4644.txt";
test_data_files[4645] = "test_data_4645.txt";
test_data_files[4646] = "test_data_4646.txt";
test_data_files[4647] = "test_data_4647.txt";
test_data_files[4648] = "test_data_4648.txt";
test_data_files[4649] = "test_data_4649.txt";
test_data_files[4650] = "test_data_4650.txt";
test_data_files[4651] = "test_data_4651.txt";
test_data_files[4652] = "test_data_4652.txt";
test_data_files[4653] = "test_data_4653.txt";
test_data_files[4654] = "test_data_4654.txt";
test_data_files[4655] = "test_data_4655.txt";
test_data_files[4656] = "test_data_4656.txt";
test_data_files[4657] = "test_data_4657.txt";
test_data_files[4658] = "test_data_4658.txt";
test_data_files[4659] = "test_data_4659.txt";
test_data_files[4660] = "test_data_4660.txt";
test_data_files[4661] = "test_data_4661.txt";
test_data_files[4662] = "test_data_4662.txt";
test_data_files[4663] = "test_data_4663.txt";
test_data_files[4664] = "test_data_4664.txt";
test_data_files[4665] = "test_data_4665.txt";
test_data_files[4666] = "test_data_4666.txt";
test_data_files[4667] = "test_data_4667.txt";
test_data_files[4668] = "test_data_4668.txt";
test_data_files[4669] = "test_data_4669.txt";
test_data_files[4670] = "test_data_4670.txt";
test_data_files[4671] = "test_data_4671.txt";
test_data_files[4672] = "test_data_4672.txt";
test_data_files[4673] = "test_data_4673.txt";
test_data_files[4674] = "test_data_4674.txt";
test_data_files[4675] = "test_data_4675.txt";
test_data_files[4676] = "test_data_4676.txt";
test_data_files[4677] = "test_data_4677.txt";
test_data_files[4678] = "test_data_4678.txt";
test_data_files[4679] = "test_data_4679.txt";
test_data_files[4680] = "test_data_4680.txt";
test_data_files[4681] = "test_data_4681.txt";
test_data_files[4682] = "test_data_4682.txt";
test_data_files[4683] = "test_data_4683.txt";
test_data_files[4684] = "test_data_4684.txt";
test_data_files[4685] = "test_data_4685.txt";
test_data_files[4686] = "test_data_4686.txt";
test_data_files[4687] = "test_data_4687.txt";
test_data_files[4688] = "test_data_4688.txt";
test_data_files[4689] = "test_data_4689.txt";
test_data_files[4690] = "test_data_4690.txt";
test_data_files[4691] = "test_data_4691.txt";
test_data_files[4692] = "test_data_4692.txt";
test_data_files[4693] = "test_data_4693.txt";
test_data_files[4694] = "test_data_4694.txt";
test_data_files[4695] = "test_data_4695.txt";
test_data_files[4696] = "test_data_4696.txt";
test_data_files[4697] = "test_data_4697.txt";
test_data_files[4698] = "test_data_4698.txt";
test_data_files[4699] = "test_data_4699.txt";
test_data_files[4700] = "test_data_4700.txt";
test_data_files[4701] = "test_data_4701.txt";
test_data_files[4702] = "test_data_4702.txt";
test_data_files[4703] = "test_data_4703.txt";
test_data_files[4704] = "test_data_4704.txt";
test_data_files[4705] = "test_data_4705.txt";
test_data_files[4706] = "test_data_4706.txt";
test_data_files[4707] = "test_data_4707.txt";
test_data_files[4708] = "test_data_4708.txt";
test_data_files[4709] = "test_data_4709.txt";
test_data_files[4710] = "test_data_4710.txt";
test_data_files[4711] = "test_data_4711.txt";
test_data_files[4712] = "test_data_4712.txt";
test_data_files[4713] = "test_data_4713.txt";
test_data_files[4714] = "test_data_4714.txt";
test_data_files[4715] = "test_data_4715.txt";
test_data_files[4716] = "test_data_4716.txt";
test_data_files[4717] = "test_data_4717.txt";
test_data_files[4718] = "test_data_4718.txt";
test_data_files[4719] = "test_data_4719.txt";
test_data_files[4720] = "test_data_4720.txt";
test_data_files[4721] = "test_data_4721.txt";
test_data_files[4722] = "test_data_4722.txt";
test_data_files[4723] = "test_data_4723.txt";
test_data_files[4724] = "test_data_4724.txt";
test_data_files[4725] = "test_data_4725.txt";
test_data_files[4726] = "test_data_4726.txt";
test_data_files[4727] = "test_data_4727.txt";
test_data_files[4728] = "test_data_4728.txt";
test_data_files[4729] = "test_data_4729.txt";
test_data_files[4730] = "test_data_4730.txt";
test_data_files[4731] = "test_data_4731.txt";
test_data_files[4732] = "test_data_4732.txt";
test_data_files[4733] = "test_data_4733.txt";
test_data_files[4734] = "test_data_4734.txt";
test_data_files[4735] = "test_data_4735.txt";
test_data_files[4736] = "test_data_4736.txt";
test_data_files[4737] = "test_data_4737.txt";
test_data_files[4738] = "test_data_4738.txt";
test_data_files[4739] = "test_data_4739.txt";
test_data_files[4740] = "test_data_4740.txt";
test_data_files[4741] = "test_data_4741.txt";
test_data_files[4742] = "test_data_4742.txt";
test_data_files[4743] = "test_data_4743.txt";
test_data_files[4744] = "test_data_4744.txt";
test_data_files[4745] = "test_data_4745.txt";
test_data_files[4746] = "test_data_4746.txt";
test_data_files[4747] = "test_data_4747.txt";
test_data_files[4748] = "test_data_4748.txt";
test_data_files[4749] = "test_data_4749.txt";
test_data_files[4750] = "test_data_4750.txt";
test_data_files[4751] = "test_data_4751.txt";
test_data_files[4752] = "test_data_4752.txt";
test_data_files[4753] = "test_data_4753.txt";
test_data_files[4754] = "test_data_4754.txt";
test_data_files[4755] = "test_data_4755.txt";
test_data_files[4756] = "test_data_4756.txt";
test_data_files[4757] = "test_data_4757.txt";
test_data_files[4758] = "test_data_4758.txt";
test_data_files[4759] = "test_data_4759.txt";
test_data_files[4760] = "test_data_4760.txt";
test_data_files[4761] = "test_data_4761.txt";
test_data_files[4762] = "test_data_4762.txt";
test_data_files[4763] = "test_data_4763.txt";
test_data_files[4764] = "test_data_4764.txt";
test_data_files[4765] = "test_data_4765.txt";
test_data_files[4766] = "test_data_4766.txt";
test_data_files[4767] = "test_data_4767.txt";
test_data_files[4768] = "test_data_4768.txt";
test_data_files[4769] = "test_data_4769.txt";
test_data_files[4770] = "test_data_4770.txt";
test_data_files[4771] = "test_data_4771.txt";
test_data_files[4772] = "test_data_4772.txt";
test_data_files[4773] = "test_data_4773.txt";
test_data_files[4774] = "test_data_4774.txt";
test_data_files[4775] = "test_data_4775.txt";
test_data_files[4776] = "test_data_4776.txt";
test_data_files[4777] = "test_data_4777.txt";
test_data_files[4778] = "test_data_4778.txt";
test_data_files[4779] = "test_data_4779.txt";
test_data_files[4780] = "test_data_4780.txt";
test_data_files[4781] = "test_data_4781.txt";
test_data_files[4782] = "test_data_4782.txt";
test_data_files[4783] = "test_data_4783.txt";
test_data_files[4784] = "test_data_4784.txt";
test_data_files[4785] = "test_data_4785.txt";
test_data_files[4786] = "test_data_4786.txt";
test_data_files[4787] = "test_data_4787.txt";
test_data_files[4788] = "test_data_4788.txt";
test_data_files[4789] = "test_data_4789.txt";
test_data_files[4790] = "test_data_4790.txt";
test_data_files[4791] = "test_data_4791.txt";
test_data_files[4792] = "test_data_4792.txt";
test_data_files[4793] = "test_data_4793.txt";
test_data_files[4794] = "test_data_4794.txt";
test_data_files[4795] = "test_data_4795.txt";
test_data_files[4796] = "test_data_4796.txt";
test_data_files[4797] = "test_data_4797.txt";
test_data_files[4798] = "test_data_4798.txt";
test_data_files[4799] = "test_data_4799.txt";
test_data_files[4800] = "test_data_4800.txt";
test_data_files[4801] = "test_data_4801.txt";
test_data_files[4802] = "test_data_4802.txt";
test_data_files[4803] = "test_data_4803.txt";
test_data_files[4804] = "test_data_4804.txt";
test_data_files[4805] = "test_data_4805.txt";
test_data_files[4806] = "test_data_4806.txt";
test_data_files[4807] = "test_data_4807.txt";
test_data_files[4808] = "test_data_4808.txt";
test_data_files[4809] = "test_data_4809.txt";
test_data_files[4810] = "test_data_4810.txt";
test_data_files[4811] = "test_data_4811.txt";
test_data_files[4812] = "test_data_4812.txt";
test_data_files[4813] = "test_data_4813.txt";
test_data_files[4814] = "test_data_4814.txt";
test_data_files[4815] = "test_data_4815.txt";
test_data_files[4816] = "test_data_4816.txt";
test_data_files[4817] = "test_data_4817.txt";
test_data_files[4818] = "test_data_4818.txt";
test_data_files[4819] = "test_data_4819.txt";
test_data_files[4820] = "test_data_4820.txt";
test_data_files[4821] = "test_data_4821.txt";
test_data_files[4822] = "test_data_4822.txt";
test_data_files[4823] = "test_data_4823.txt";
test_data_files[4824] = "test_data_4824.txt";
test_data_files[4825] = "test_data_4825.txt";
test_data_files[4826] = "test_data_4826.txt";
test_data_files[4827] = "test_data_4827.txt";
test_data_files[4828] = "test_data_4828.txt";
test_data_files[4829] = "test_data_4829.txt";
test_data_files[4830] = "test_data_4830.txt";
test_data_files[4831] = "test_data_4831.txt";
test_data_files[4832] = "test_data_4832.txt";
test_data_files[4833] = "test_data_4833.txt";
test_data_files[4834] = "test_data_4834.txt";
test_data_files[4835] = "test_data_4835.txt";
test_data_files[4836] = "test_data_4836.txt";
test_data_files[4837] = "test_data_4837.txt";
test_data_files[4838] = "test_data_4838.txt";
test_data_files[4839] = "test_data_4839.txt";
test_data_files[4840] = "test_data_4840.txt";
test_data_files[4841] = "test_data_4841.txt";
test_data_files[4842] = "test_data_4842.txt";
test_data_files[4843] = "test_data_4843.txt";
test_data_files[4844] = "test_data_4844.txt";
test_data_files[4845] = "test_data_4845.txt";
test_data_files[4846] = "test_data_4846.txt";
test_data_files[4847] = "test_data_4847.txt";
test_data_files[4848] = "test_data_4848.txt";
test_data_files[4849] = "test_data_4849.txt";
test_data_files[4850] = "test_data_4850.txt";
test_data_files[4851] = "test_data_4851.txt";
test_data_files[4852] = "test_data_4852.txt";
test_data_files[4853] = "test_data_4853.txt";
test_data_files[4854] = "test_data_4854.txt";
test_data_files[4855] = "test_data_4855.txt";
test_data_files[4856] = "test_data_4856.txt";
test_data_files[4857] = "test_data_4857.txt";
test_data_files[4858] = "test_data_4858.txt";
test_data_files[4859] = "test_data_4859.txt";
test_data_files[4860] = "test_data_4860.txt";
test_data_files[4861] = "test_data_4861.txt";
test_data_files[4862] = "test_data_4862.txt";
test_data_files[4863] = "test_data_4863.txt";
test_data_files[4864] = "test_data_4864.txt";
test_data_files[4865] = "test_data_4865.txt";
test_data_files[4866] = "test_data_4866.txt";
test_data_files[4867] = "test_data_4867.txt";
test_data_files[4868] = "test_data_4868.txt";
test_data_files[4869] = "test_data_4869.txt";
test_data_files[4870] = "test_data_4870.txt";
test_data_files[4871] = "test_data_4871.txt";
test_data_files[4872] = "test_data_4872.txt";
test_data_files[4873] = "test_data_4873.txt";
test_data_files[4874] = "test_data_4874.txt";
test_data_files[4875] = "test_data_4875.txt";
test_data_files[4876] = "test_data_4876.txt";
test_data_files[4877] = "test_data_4877.txt";
test_data_files[4878] = "test_data_4878.txt";
test_data_files[4879] = "test_data_4879.txt";
test_data_files[4880] = "test_data_4880.txt";
test_data_files[4881] = "test_data_4881.txt";
test_data_files[4882] = "test_data_4882.txt";
test_data_files[4883] = "test_data_4883.txt";
test_data_files[4884] = "test_data_4884.txt";
test_data_files[4885] = "test_data_4885.txt";
test_data_files[4886] = "test_data_4886.txt";
test_data_files[4887] = "test_data_4887.txt";
test_data_files[4888] = "test_data_4888.txt";
test_data_files[4889] = "test_data_4889.txt";
test_data_files[4890] = "test_data_4890.txt";
test_data_files[4891] = "test_data_4891.txt";
test_data_files[4892] = "test_data_4892.txt";
test_data_files[4893] = "test_data_4893.txt";
test_data_files[4894] = "test_data_4894.txt";
test_data_files[4895] = "test_data_4895.txt";
test_data_files[4896] = "test_data_4896.txt";
test_data_files[4897] = "test_data_4897.txt";
test_data_files[4898] = "test_data_4898.txt";
test_data_files[4899] = "test_data_4899.txt";
test_data_files[4900] = "test_data_4900.txt";
test_data_files[4901] = "test_data_4901.txt";
test_data_files[4902] = "test_data_4902.txt";
test_data_files[4903] = "test_data_4903.txt";
test_data_files[4904] = "test_data_4904.txt";
test_data_files[4905] = "test_data_4905.txt";
test_data_files[4906] = "test_data_4906.txt";
test_data_files[4907] = "test_data_4907.txt";
test_data_files[4908] = "test_data_4908.txt";
test_data_files[4909] = "test_data_4909.txt";
test_data_files[4910] = "test_data_4910.txt";
test_data_files[4911] = "test_data_4911.txt";
test_data_files[4912] = "test_data_4912.txt";
test_data_files[4913] = "test_data_4913.txt";
test_data_files[4914] = "test_data_4914.txt";
test_data_files[4915] = "test_data_4915.txt";
test_data_files[4916] = "test_data_4916.txt";
test_data_files[4917] = "test_data_4917.txt";
test_data_files[4918] = "test_data_4918.txt";
test_data_files[4919] = "test_data_4919.txt";
test_data_files[4920] = "test_data_4920.txt";
test_data_files[4921] = "test_data_4921.txt";
test_data_files[4922] = "test_data_4922.txt";
test_data_files[4923] = "test_data_4923.txt";
test_data_files[4924] = "test_data_4924.txt";
test_data_files[4925] = "test_data_4925.txt";
test_data_files[4926] = "test_data_4926.txt";
test_data_files[4927] = "test_data_4927.txt";
test_data_files[4928] = "test_data_4928.txt";
test_data_files[4929] = "test_data_4929.txt";
test_data_files[4930] = "test_data_4930.txt";
test_data_files[4931] = "test_data_4931.txt";
test_data_files[4932] = "test_data_4932.txt";
test_data_files[4933] = "test_data_4933.txt";
test_data_files[4934] = "test_data_4934.txt";
test_data_files[4935] = "test_data_4935.txt";
test_data_files[4936] = "test_data_4936.txt";
test_data_files[4937] = "test_data_4937.txt";
test_data_files[4938] = "test_data_4938.txt";
test_data_files[4939] = "test_data_4939.txt";
test_data_files[4940] = "test_data_4940.txt";
test_data_files[4941] = "test_data_4941.txt";
test_data_files[4942] = "test_data_4942.txt";
test_data_files[4943] = "test_data_4943.txt";
test_data_files[4944] = "test_data_4944.txt";
test_data_files[4945] = "test_data_4945.txt";
test_data_files[4946] = "test_data_4946.txt";
test_data_files[4947] = "test_data_4947.txt";
test_data_files[4948] = "test_data_4948.txt";
test_data_files[4949] = "test_data_4949.txt";
test_data_files[4950] = "test_data_4950.txt";
test_data_files[4951] = "test_data_4951.txt";
test_data_files[4952] = "test_data_4952.txt";
test_data_files[4953] = "test_data_4953.txt";
test_data_files[4954] = "test_data_4954.txt";
test_data_files[4955] = "test_data_4955.txt";
test_data_files[4956] = "test_data_4956.txt";
test_data_files[4957] = "test_data_4957.txt";
test_data_files[4958] = "test_data_4958.txt";
test_data_files[4959] = "test_data_4959.txt";
test_data_files[4960] = "test_data_4960.txt";
test_data_files[4961] = "test_data_4961.txt";
test_data_files[4962] = "test_data_4962.txt";
test_data_files[4963] = "test_data_4963.txt";
test_data_files[4964] = "test_data_4964.txt";
test_data_files[4965] = "test_data_4965.txt";
test_data_files[4966] = "test_data_4966.txt";
test_data_files[4967] = "test_data_4967.txt";
test_data_files[4968] = "test_data_4968.txt";
test_data_files[4969] = "test_data_4969.txt";
test_data_files[4970] = "test_data_4970.txt";
test_data_files[4971] = "test_data_4971.txt";
test_data_files[4972] = "test_data_4972.txt";
test_data_files[4973] = "test_data_4973.txt";
test_data_files[4974] = "test_data_4974.txt";
test_data_files[4975] = "test_data_4975.txt";
test_data_files[4976] = "test_data_4976.txt";
test_data_files[4977] = "test_data_4977.txt";
test_data_files[4978] = "test_data_4978.txt";
test_data_files[4979] = "test_data_4979.txt";
test_data_files[4980] = "test_data_4980.txt";
test_data_files[4981] = "test_data_4981.txt";
test_data_files[4982] = "test_data_4982.txt";
test_data_files[4983] = "test_data_4983.txt";
test_data_files[4984] = "test_data_4984.txt";
test_data_files[4985] = "test_data_4985.txt";
test_data_files[4986] = "test_data_4986.txt";
test_data_files[4987] = "test_data_4987.txt";
test_data_files[4988] = "test_data_4988.txt";
test_data_files[4989] = "test_data_4989.txt";
test_data_files[4990] = "test_data_4990.txt";
test_data_files[4991] = "test_data_4991.txt";
test_data_files[4992] = "test_data_4992.txt";
test_data_files[4993] = "test_data_4993.txt";
test_data_files[4994] = "test_data_4994.txt";
test_data_files[4995] = "test_data_4995.txt";
test_data_files[4996] = "test_data_4996.txt";
test_data_files[4997] = "test_data_4997.txt";
test_data_files[4998] = "test_data_4998.txt";
test_data_files[4999] = "test_data_4999.txt";
test_data_files[5000] = "test_data_5000.txt";
test_data_files[5001] = "test_data_5001.txt";
test_data_files[5002] = "test_data_5002.txt";
test_data_files[5003] = "test_data_5003.txt";
test_data_files[5004] = "test_data_5004.txt";
test_data_files[5005] = "test_data_5005.txt";
test_data_files[5006] = "test_data_5006.txt";
test_data_files[5007] = "test_data_5007.txt";
test_data_files[5008] = "test_data_5008.txt";
test_data_files[5009] = "test_data_5009.txt";
test_data_files[5010] = "test_data_5010.txt";
test_data_files[5011] = "test_data_5011.txt";
test_data_files[5012] = "test_data_5012.txt";
test_data_files[5013] = "test_data_5013.txt";
test_data_files[5014] = "test_data_5014.txt";
test_data_files[5015] = "test_data_5015.txt";
test_data_files[5016] = "test_data_5016.txt";
test_data_files[5017] = "test_data_5017.txt";
test_data_files[5018] = "test_data_5018.txt";
test_data_files[5019] = "test_data_5019.txt";
test_data_files[5020] = "test_data_5020.txt";
test_data_files[5021] = "test_data_5021.txt";
test_data_files[5022] = "test_data_5022.txt";
test_data_files[5023] = "test_data_5023.txt";
test_data_files[5024] = "test_data_5024.txt";
test_data_files[5025] = "test_data_5025.txt";
test_data_files[5026] = "test_data_5026.txt";
test_data_files[5027] = "test_data_5027.txt";
test_data_files[5028] = "test_data_5028.txt";
test_data_files[5029] = "test_data_5029.txt";
test_data_files[5030] = "test_data_5030.txt";
test_data_files[5031] = "test_data_5031.txt";
test_data_files[5032] = "test_data_5032.txt";
test_data_files[5033] = "test_data_5033.txt";
test_data_files[5034] = "test_data_5034.txt";
test_data_files[5035] = "test_data_5035.txt";
test_data_files[5036] = "test_data_5036.txt";
test_data_files[5037] = "test_data_5037.txt";
test_data_files[5038] = "test_data_5038.txt";
test_data_files[5039] = "test_data_5039.txt";
test_data_files[5040] = "test_data_5040.txt";
test_data_files[5041] = "test_data_5041.txt";
test_data_files[5042] = "test_data_5042.txt";
test_data_files[5043] = "test_data_5043.txt";
test_data_files[5044] = "test_data_5044.txt";
test_data_files[5045] = "test_data_5045.txt";
test_data_files[5046] = "test_data_5046.txt";
test_data_files[5047] = "test_data_5047.txt";
test_data_files[5048] = "test_data_5048.txt";
test_data_files[5049] = "test_data_5049.txt";
test_data_files[5050] = "test_data_5050.txt";
test_data_files[5051] = "test_data_5051.txt";
test_data_files[5052] = "test_data_5052.txt";
test_data_files[5053] = "test_data_5053.txt";
test_data_files[5054] = "test_data_5054.txt";
test_data_files[5055] = "test_data_5055.txt";
test_data_files[5056] = "test_data_5056.txt";
test_data_files[5057] = "test_data_5057.txt";
test_data_files[5058] = "test_data_5058.txt";
test_data_files[5059] = "test_data_5059.txt";
test_data_files[5060] = "test_data_5060.txt";
test_data_files[5061] = "test_data_5061.txt";
test_data_files[5062] = "test_data_5062.txt";
test_data_files[5063] = "test_data_5063.txt";
test_data_files[5064] = "test_data_5064.txt";
test_data_files[5065] = "test_data_5065.txt";
test_data_files[5066] = "test_data_5066.txt";
test_data_files[5067] = "test_data_5067.txt";
test_data_files[5068] = "test_data_5068.txt";
test_data_files[5069] = "test_data_5069.txt";
test_data_files[5070] = "test_data_5070.txt";
test_data_files[5071] = "test_data_5071.txt";
test_data_files[5072] = "test_data_5072.txt";
test_data_files[5073] = "test_data_5073.txt";
test_data_files[5074] = "test_data_5074.txt";
test_data_files[5075] = "test_data_5075.txt";
test_data_files[5076] = "test_data_5076.txt";
test_data_files[5077] = "test_data_5077.txt";
test_data_files[5078] = "test_data_5078.txt";
test_data_files[5079] = "test_data_5079.txt";
test_data_files[5080] = "test_data_5080.txt";
test_data_files[5081] = "test_data_5081.txt";
test_data_files[5082] = "test_data_5082.txt";
test_data_files[5083] = "test_data_5083.txt";
test_data_files[5084] = "test_data_5084.txt";
test_data_files[5085] = "test_data_5085.txt";
test_data_files[5086] = "test_data_5086.txt";
test_data_files[5087] = "test_data_5087.txt";
test_data_files[5088] = "test_data_5088.txt";
test_data_files[5089] = "test_data_5089.txt";
test_data_files[5090] = "test_data_5090.txt";
test_data_files[5091] = "test_data_5091.txt";
test_data_files[5092] = "test_data_5092.txt";
test_data_files[5093] = "test_data_5093.txt";
test_data_files[5094] = "test_data_5094.txt";
test_data_files[5095] = "test_data_5095.txt";
test_data_files[5096] = "test_data_5096.txt";
test_data_files[5097] = "test_data_5097.txt";
test_data_files[5098] = "test_data_5098.txt";
test_data_files[5099] = "test_data_5099.txt";
test_data_files[5100] = "test_data_5100.txt";
test_data_files[5101] = "test_data_5101.txt";
test_data_files[5102] = "test_data_5102.txt";
test_data_files[5103] = "test_data_5103.txt";
test_data_files[5104] = "test_data_5104.txt";
test_data_files[5105] = "test_data_5105.txt";
test_data_files[5106] = "test_data_5106.txt";
test_data_files[5107] = "test_data_5107.txt";
test_data_files[5108] = "test_data_5108.txt";
test_data_files[5109] = "test_data_5109.txt";
test_data_files[5110] = "test_data_5110.txt";
test_data_files[5111] = "test_data_5111.txt";
test_data_files[5112] = "test_data_5112.txt";
test_data_files[5113] = "test_data_5113.txt";
test_data_files[5114] = "test_data_5114.txt";
test_data_files[5115] = "test_data_5115.txt";
test_data_files[5116] = "test_data_5116.txt";
test_data_files[5117] = "test_data_5117.txt";
test_data_files[5118] = "test_data_5118.txt";
test_data_files[5119] = "test_data_5119.txt";
test_data_files[5120] = "test_data_5120.txt";
test_data_files[5121] = "test_data_5121.txt";
test_data_files[5122] = "test_data_5122.txt";
test_data_files[5123] = "test_data_5123.txt";
test_data_files[5124] = "test_data_5124.txt";
test_data_files[5125] = "test_data_5125.txt";
test_data_files[5126] = "test_data_5126.txt";
test_data_files[5127] = "test_data_5127.txt";
test_data_files[5128] = "test_data_5128.txt";
test_data_files[5129] = "test_data_5129.txt";
test_data_files[5130] = "test_data_5130.txt";
test_data_files[5131] = "test_data_5131.txt";
test_data_files[5132] = "test_data_5132.txt";
test_data_files[5133] = "test_data_5133.txt";
test_data_files[5134] = "test_data_5134.txt";
test_data_files[5135] = "test_data_5135.txt";
test_data_files[5136] = "test_data_5136.txt";
test_data_files[5137] = "test_data_5137.txt";
test_data_files[5138] = "test_data_5138.txt";
test_data_files[5139] = "test_data_5139.txt";
test_data_files[5140] = "test_data_5140.txt";
test_data_files[5141] = "test_data_5141.txt";
test_data_files[5142] = "test_data_5142.txt";
test_data_files[5143] = "test_data_5143.txt";
test_data_files[5144] = "test_data_5144.txt";
test_data_files[5145] = "test_data_5145.txt";
test_data_files[5146] = "test_data_5146.txt";
test_data_files[5147] = "test_data_5147.txt";
test_data_files[5148] = "test_data_5148.txt";
test_data_files[5149] = "test_data_5149.txt";
test_data_files[5150] = "test_data_5150.txt";
test_data_files[5151] = "test_data_5151.txt";
test_data_files[5152] = "test_data_5152.txt";
test_data_files[5153] = "test_data_5153.txt";
test_data_files[5154] = "test_data_5154.txt";
test_data_files[5155] = "test_data_5155.txt";
test_data_files[5156] = "test_data_5156.txt";
test_data_files[5157] = "test_data_5157.txt";
test_data_files[5158] = "test_data_5158.txt";
test_data_files[5159] = "test_data_5159.txt";
test_data_files[5160] = "test_data_5160.txt";
test_data_files[5161] = "test_data_5161.txt";
test_data_files[5162] = "test_data_5162.txt";
test_data_files[5163] = "test_data_5163.txt";
test_data_files[5164] = "test_data_5164.txt";
test_data_files[5165] = "test_data_5165.txt";
test_data_files[5166] = "test_data_5166.txt";
test_data_files[5167] = "test_data_5167.txt";
test_data_files[5168] = "test_data_5168.txt";
test_data_files[5169] = "test_data_5169.txt";
test_data_files[5170] = "test_data_5170.txt";
test_data_files[5171] = "test_data_5171.txt";
test_data_files[5172] = "test_data_5172.txt";
test_data_files[5173] = "test_data_5173.txt";
test_data_files[5174] = "test_data_5174.txt";
test_data_files[5175] = "test_data_5175.txt";
test_data_files[5176] = "test_data_5176.txt";
test_data_files[5177] = "test_data_5177.txt";
test_data_files[5178] = "test_data_5178.txt";
test_data_files[5179] = "test_data_5179.txt";
test_data_files[5180] = "test_data_5180.txt";
test_data_files[5181] = "test_data_5181.txt";
test_data_files[5182] = "test_data_5182.txt";
test_data_files[5183] = "test_data_5183.txt";
test_data_files[5184] = "test_data_5184.txt";
test_data_files[5185] = "test_data_5185.txt";
test_data_files[5186] = "test_data_5186.txt";
test_data_files[5187] = "test_data_5187.txt";
test_data_files[5188] = "test_data_5188.txt";
test_data_files[5189] = "test_data_5189.txt";
test_data_files[5190] = "test_data_5190.txt";
test_data_files[5191] = "test_data_5191.txt";
test_data_files[5192] = "test_data_5192.txt";
test_data_files[5193] = "test_data_5193.txt";
test_data_files[5194] = "test_data_5194.txt";
test_data_files[5195] = "test_data_5195.txt";
test_data_files[5196] = "test_data_5196.txt";
test_data_files[5197] = "test_data_5197.txt";
test_data_files[5198] = "test_data_5198.txt";
test_data_files[5199] = "test_data_5199.txt";
test_data_files[5200] = "test_data_5200.txt";
test_data_files[5201] = "test_data_5201.txt";
test_data_files[5202] = "test_data_5202.txt";
test_data_files[5203] = "test_data_5203.txt";
test_data_files[5204] = "test_data_5204.txt";
test_data_files[5205] = "test_data_5205.txt";
test_data_files[5206] = "test_data_5206.txt";
test_data_files[5207] = "test_data_5207.txt";
test_data_files[5208] = "test_data_5208.txt";
test_data_files[5209] = "test_data_5209.txt";
test_data_files[5210] = "test_data_5210.txt";
test_data_files[5211] = "test_data_5211.txt";
test_data_files[5212] = "test_data_5212.txt";
test_data_files[5213] = "test_data_5213.txt";
test_data_files[5214] = "test_data_5214.txt";
test_data_files[5215] = "test_data_5215.txt";
test_data_files[5216] = "test_data_5216.txt";
test_data_files[5217] = "test_data_5217.txt";
test_data_files[5218] = "test_data_5218.txt";
test_data_files[5219] = "test_data_5219.txt";
test_data_files[5220] = "test_data_5220.txt";
test_data_files[5221] = "test_data_5221.txt";
test_data_files[5222] = "test_data_5222.txt";
test_data_files[5223] = "test_data_5223.txt";
test_data_files[5224] = "test_data_5224.txt";
test_data_files[5225] = "test_data_5225.txt";
test_data_files[5226] = "test_data_5226.txt";
test_data_files[5227] = "test_data_5227.txt";
test_data_files[5228] = "test_data_5228.txt";
test_data_files[5229] = "test_data_5229.txt";
test_data_files[5230] = "test_data_5230.txt";
test_data_files[5231] = "test_data_5231.txt";
test_data_files[5232] = "test_data_5232.txt";
test_data_files[5233] = "test_data_5233.txt";
test_data_files[5234] = "test_data_5234.txt";
test_data_files[5235] = "test_data_5235.txt";
test_data_files[5236] = "test_data_5236.txt";
test_data_files[5237] = "test_data_5237.txt";
test_data_files[5238] = "test_data_5238.txt";
test_data_files[5239] = "test_data_5239.txt";
test_data_files[5240] = "test_data_5240.txt";
test_data_files[5241] = "test_data_5241.txt";
test_data_files[5242] = "test_data_5242.txt";
test_data_files[5243] = "test_data_5243.txt";
test_data_files[5244] = "test_data_5244.txt";
test_data_files[5245] = "test_data_5245.txt";
test_data_files[5246] = "test_data_5246.txt";
test_data_files[5247] = "test_data_5247.txt";
test_data_files[5248] = "test_data_5248.txt";
test_data_files[5249] = "test_data_5249.txt";
test_data_files[5250] = "test_data_5250.txt";
test_data_files[5251] = "test_data_5251.txt";
test_data_files[5252] = "test_data_5252.txt";
test_data_files[5253] = "test_data_5253.txt";
test_data_files[5254] = "test_data_5254.txt";
test_data_files[5255] = "test_data_5255.txt";
test_data_files[5256] = "test_data_5256.txt";
test_data_files[5257] = "test_data_5257.txt";
test_data_files[5258] = "test_data_5258.txt";
test_data_files[5259] = "test_data_5259.txt";
test_data_files[5260] = "test_data_5260.txt";
test_data_files[5261] = "test_data_5261.txt";
test_data_files[5262] = "test_data_5262.txt";
test_data_files[5263] = "test_data_5263.txt";
test_data_files[5264] = "test_data_5264.txt";
test_data_files[5265] = "test_data_5265.txt";
test_data_files[5266] = "test_data_5266.txt";
test_data_files[5267] = "test_data_5267.txt";
test_data_files[5268] = "test_data_5268.txt";
test_data_files[5269] = "test_data_5269.txt";
test_data_files[5270] = "test_data_5270.txt";
test_data_files[5271] = "test_data_5271.txt";
test_data_files[5272] = "test_data_5272.txt";
test_data_files[5273] = "test_data_5273.txt";
test_data_files[5274] = "test_data_5274.txt";
test_data_files[5275] = "test_data_5275.txt";
test_data_files[5276] = "test_data_5276.txt";
test_data_files[5277] = "test_data_5277.txt";
test_data_files[5278] = "test_data_5278.txt";
test_data_files[5279] = "test_data_5279.txt";
test_data_files[5280] = "test_data_5280.txt";
test_data_files[5281] = "test_data_5281.txt";
test_data_files[5282] = "test_data_5282.txt";
test_data_files[5283] = "test_data_5283.txt";
test_data_files[5284] = "test_data_5284.txt";
test_data_files[5285] = "test_data_5285.txt";
test_data_files[5286] = "test_data_5286.txt";
test_data_files[5287] = "test_data_5287.txt";
test_data_files[5288] = "test_data_5288.txt";
test_data_files[5289] = "test_data_5289.txt";
test_data_files[5290] = "test_data_5290.txt";
test_data_files[5291] = "test_data_5291.txt";
test_data_files[5292] = "test_data_5292.txt";
test_data_files[5293] = "test_data_5293.txt";
test_data_files[5294] = "test_data_5294.txt";
test_data_files[5295] = "test_data_5295.txt";
test_data_files[5296] = "test_data_5296.txt";
test_data_files[5297] = "test_data_5297.txt";
test_data_files[5298] = "test_data_5298.txt";
test_data_files[5299] = "test_data_5299.txt";
test_data_files[5300] = "test_data_5300.txt";
test_data_files[5301] = "test_data_5301.txt";
test_data_files[5302] = "test_data_5302.txt";
test_data_files[5303] = "test_data_5303.txt";
test_data_files[5304] = "test_data_5304.txt";
test_data_files[5305] = "test_data_5305.txt";
test_data_files[5306] = "test_data_5306.txt";
test_data_files[5307] = "test_data_5307.txt";
test_data_files[5308] = "test_data_5308.txt";
test_data_files[5309] = "test_data_5309.txt";
test_data_files[5310] = "test_data_5310.txt";
test_data_files[5311] = "test_data_5311.txt";
test_data_files[5312] = "test_data_5312.txt";
test_data_files[5313] = "test_data_5313.txt";
test_data_files[5314] = "test_data_5314.txt";
test_data_files[5315] = "test_data_5315.txt";
test_data_files[5316] = "test_data_5316.txt";
test_data_files[5317] = "test_data_5317.txt";
test_data_files[5318] = "test_data_5318.txt";
test_data_files[5319] = "test_data_5319.txt";
test_data_files[5320] = "test_data_5320.txt";
test_data_files[5321] = "test_data_5321.txt";
test_data_files[5322] = "test_data_5322.txt";
test_data_files[5323] = "test_data_5323.txt";
test_data_files[5324] = "test_data_5324.txt";
test_data_files[5325] = "test_data_5325.txt";
test_data_files[5326] = "test_data_5326.txt";
test_data_files[5327] = "test_data_5327.txt";
test_data_files[5328] = "test_data_5328.txt";
test_data_files[5329] = "test_data_5329.txt";
test_data_files[5330] = "test_data_5330.txt";
test_data_files[5331] = "test_data_5331.txt";
test_data_files[5332] = "test_data_5332.txt";
test_data_files[5333] = "test_data_5333.txt";
test_data_files[5334] = "test_data_5334.txt";
test_data_files[5335] = "test_data_5335.txt";
test_data_files[5336] = "test_data_5336.txt";
test_data_files[5337] = "test_data_5337.txt";
test_data_files[5338] = "test_data_5338.txt";
test_data_files[5339] = "test_data_5339.txt";
test_data_files[5340] = "test_data_5340.txt";
test_data_files[5341] = "test_data_5341.txt";
test_data_files[5342] = "test_data_5342.txt";
test_data_files[5343] = "test_data_5343.txt";
test_data_files[5344] = "test_data_5344.txt";
test_data_files[5345] = "test_data_5345.txt";
test_data_files[5346] = "test_data_5346.txt";
test_data_files[5347] = "test_data_5347.txt";
test_data_files[5348] = "test_data_5348.txt";
test_data_files[5349] = "test_data_5349.txt";
test_data_files[5350] = "test_data_5350.txt";
test_data_files[5351] = "test_data_5351.txt";
test_data_files[5352] = "test_data_5352.txt";
test_data_files[5353] = "test_data_5353.txt";
test_data_files[5354] = "test_data_5354.txt";
test_data_files[5355] = "test_data_5355.txt";
test_data_files[5356] = "test_data_5356.txt";
test_data_files[5357] = "test_data_5357.txt";
test_data_files[5358] = "test_data_5358.txt";
test_data_files[5359] = "test_data_5359.txt";
test_data_files[5360] = "test_data_5360.txt";
test_data_files[5361] = "test_data_5361.txt";
test_data_files[5362] = "test_data_5362.txt";
test_data_files[5363] = "test_data_5363.txt";
test_data_files[5364] = "test_data_5364.txt";
test_data_files[5365] = "test_data_5365.txt";
test_data_files[5366] = "test_data_5366.txt";
test_data_files[5367] = "test_data_5367.txt";
test_data_files[5368] = "test_data_5368.txt";
test_data_files[5369] = "test_data_5369.txt";
test_data_files[5370] = "test_data_5370.txt";
test_data_files[5371] = "test_data_5371.txt";
test_data_files[5372] = "test_data_5372.txt";
test_data_files[5373] = "test_data_5373.txt";
test_data_files[5374] = "test_data_5374.txt";
test_data_files[5375] = "test_data_5375.txt";
test_data_files[5376] = "test_data_5376.txt";
test_data_files[5377] = "test_data_5377.txt";
test_data_files[5378] = "test_data_5378.txt";
test_data_files[5379] = "test_data_5379.txt";
test_data_files[5380] = "test_data_5380.txt";
test_data_files[5381] = "test_data_5381.txt";
test_data_files[5382] = "test_data_5382.txt";
test_data_files[5383] = "test_data_5383.txt";
test_data_files[5384] = "test_data_5384.txt";
test_data_files[5385] = "test_data_5385.txt";
test_data_files[5386] = "test_data_5386.txt";
test_data_files[5387] = "test_data_5387.txt";
test_data_files[5388] = "test_data_5388.txt";
test_data_files[5389] = "test_data_5389.txt";
test_data_files[5390] = "test_data_5390.txt";
test_data_files[5391] = "test_data_5391.txt";
test_data_files[5392] = "test_data_5392.txt";
test_data_files[5393] = "test_data_5393.txt";
test_data_files[5394] = "test_data_5394.txt";
test_data_files[5395] = "test_data_5395.txt";
test_data_files[5396] = "test_data_5396.txt";
test_data_files[5397] = "test_data_5397.txt";
test_data_files[5398] = "test_data_5398.txt";
test_data_files[5399] = "test_data_5399.txt";
test_data_files[5400] = "test_data_5400.txt";
test_data_files[5401] = "test_data_5401.txt";
test_data_files[5402] = "test_data_5402.txt";
test_data_files[5403] = "test_data_5403.txt";
test_data_files[5404] = "test_data_5404.txt";
test_data_files[5405] = "test_data_5405.txt";
test_data_files[5406] = "test_data_5406.txt";
test_data_files[5407] = "test_data_5407.txt";
test_data_files[5408] = "test_data_5408.txt";
test_data_files[5409] = "test_data_5409.txt";
test_data_files[5410] = "test_data_5410.txt";
test_data_files[5411] = "test_data_5411.txt";
test_data_files[5412] = "test_data_5412.txt";
test_data_files[5413] = "test_data_5413.txt";
test_data_files[5414] = "test_data_5414.txt";
test_data_files[5415] = "test_data_5415.txt";
test_data_files[5416] = "test_data_5416.txt";
test_data_files[5417] = "test_data_5417.txt";
test_data_files[5418] = "test_data_5418.txt";
test_data_files[5419] = "test_data_5419.txt";
test_data_files[5420] = "test_data_5420.txt";
test_data_files[5421] = "test_data_5421.txt";
test_data_files[5422] = "test_data_5422.txt";
test_data_files[5423] = "test_data_5423.txt";
test_data_files[5424] = "test_data_5424.txt";
test_data_files[5425] = "test_data_5425.txt";
test_data_files[5426] = "test_data_5426.txt";
test_data_files[5427] = "test_data_5427.txt";
test_data_files[5428] = "test_data_5428.txt";
test_data_files[5429] = "test_data_5429.txt";
test_data_files[5430] = "test_data_5430.txt";
test_data_files[5431] = "test_data_5431.txt";
test_data_files[5432] = "test_data_5432.txt";
test_data_files[5433] = "test_data_5433.txt";
test_data_files[5434] = "test_data_5434.txt";
test_data_files[5435] = "test_data_5435.txt";
test_data_files[5436] = "test_data_5436.txt";
test_data_files[5437] = "test_data_5437.txt";
test_data_files[5438] = "test_data_5438.txt";
test_data_files[5439] = "test_data_5439.txt";
test_data_files[5440] = "test_data_5440.txt";
test_data_files[5441] = "test_data_5441.txt";
test_data_files[5442] = "test_data_5442.txt";
test_data_files[5443] = "test_data_5443.txt";
test_data_files[5444] = "test_data_5444.txt";
test_data_files[5445] = "test_data_5445.txt";
test_data_files[5446] = "test_data_5446.txt";
test_data_files[5447] = "test_data_5447.txt";
test_data_files[5448] = "test_data_5448.txt";
test_data_files[5449] = "test_data_5449.txt";
test_data_files[5450] = "test_data_5450.txt";
test_data_files[5451] = "test_data_5451.txt";
test_data_files[5452] = "test_data_5452.txt";
test_data_files[5453] = "test_data_5453.txt";
test_data_files[5454] = "test_data_5454.txt";
test_data_files[5455] = "test_data_5455.txt";
test_data_files[5456] = "test_data_5456.txt";
test_data_files[5457] = "test_data_5457.txt";
test_data_files[5458] = "test_data_5458.txt";
test_data_files[5459] = "test_data_5459.txt";
test_data_files[5460] = "test_data_5460.txt";
test_data_files[5461] = "test_data_5461.txt";
test_data_files[5462] = "test_data_5462.txt";
test_data_files[5463] = "test_data_5463.txt";
test_data_files[5464] = "test_data_5464.txt";
test_data_files[5465] = "test_data_5465.txt";
test_data_files[5466] = "test_data_5466.txt";
test_data_files[5467] = "test_data_5467.txt";
test_data_files[5468] = "test_data_5468.txt";
test_data_files[5469] = "test_data_5469.txt";
test_data_files[5470] = "test_data_5470.txt";
test_data_files[5471] = "test_data_5471.txt";
test_data_files[5472] = "test_data_5472.txt";
test_data_files[5473] = "test_data_5473.txt";
test_data_files[5474] = "test_data_5474.txt";
test_data_files[5475] = "test_data_5475.txt";
test_data_files[5476] = "test_data_5476.txt";
test_data_files[5477] = "test_data_5477.txt";
test_data_files[5478] = "test_data_5478.txt";
test_data_files[5479] = "test_data_5479.txt";
test_data_files[5480] = "test_data_5480.txt";
test_data_files[5481] = "test_data_5481.txt";
test_data_files[5482] = "test_data_5482.txt";
test_data_files[5483] = "test_data_5483.txt";
test_data_files[5484] = "test_data_5484.txt";
test_data_files[5485] = "test_data_5485.txt";
test_data_files[5486] = "test_data_5486.txt";
test_data_files[5487] = "test_data_5487.txt";
test_data_files[5488] = "test_data_5488.txt";
test_data_files[5489] = "test_data_5489.txt";
test_data_files[5490] = "test_data_5490.txt";
test_data_files[5491] = "test_data_5491.txt";
test_data_files[5492] = "test_data_5492.txt";
test_data_files[5493] = "test_data_5493.txt";
test_data_files[5494] = "test_data_5494.txt";
test_data_files[5495] = "test_data_5495.txt";
test_data_files[5496] = "test_data_5496.txt";
test_data_files[5497] = "test_data_5497.txt";
test_data_files[5498] = "test_data_5498.txt";
test_data_files[5499] = "test_data_5499.txt";
test_data_files[5500] = "test_data_5500.txt";
test_data_files[5501] = "test_data_5501.txt";
test_data_files[5502] = "test_data_5502.txt";
test_data_files[5503] = "test_data_5503.txt";
test_data_files[5504] = "test_data_5504.txt";
test_data_files[5505] = "test_data_5505.txt";
test_data_files[5506] = "test_data_5506.txt";
test_data_files[5507] = "test_data_5507.txt";
test_data_files[5508] = "test_data_5508.txt";
test_data_files[5509] = "test_data_5509.txt";
test_data_files[5510] = "test_data_5510.txt";
test_data_files[5511] = "test_data_5511.txt";
test_data_files[5512] = "test_data_5512.txt";
test_data_files[5513] = "test_data_5513.txt";
test_data_files[5514] = "test_data_5514.txt";
test_data_files[5515] = "test_data_5515.txt";
test_data_files[5516] = "test_data_5516.txt";
test_data_files[5517] = "test_data_5517.txt";
test_data_files[5518] = "test_data_5518.txt";
test_data_files[5519] = "test_data_5519.txt";
test_data_files[5520] = "test_data_5520.txt";
test_data_files[5521] = "test_data_5521.txt";
test_data_files[5522] = "test_data_5522.txt";
test_data_files[5523] = "test_data_5523.txt";
test_data_files[5524] = "test_data_5524.txt";
test_data_files[5525] = "test_data_5525.txt";
test_data_files[5526] = "test_data_5526.txt";
test_data_files[5527] = "test_data_5527.txt";
test_data_files[5528] = "test_data_5528.txt";
test_data_files[5529] = "test_data_5529.txt";
test_data_files[5530] = "test_data_5530.txt";
test_data_files[5531] = "test_data_5531.txt";
test_data_files[5532] = "test_data_5532.txt";
test_data_files[5533] = "test_data_5533.txt";
test_data_files[5534] = "test_data_5534.txt";
test_data_files[5535] = "test_data_5535.txt";
test_data_files[5536] = "test_data_5536.txt";
test_data_files[5537] = "test_data_5537.txt";
test_data_files[5538] = "test_data_5538.txt";
test_data_files[5539] = "test_data_5539.txt";
test_data_files[5540] = "test_data_5540.txt";
test_data_files[5541] = "test_data_5541.txt";
test_data_files[5542] = "test_data_5542.txt";
test_data_files[5543] = "test_data_5543.txt";
test_data_files[5544] = "test_data_5544.txt";
test_data_files[5545] = "test_data_5545.txt";
test_data_files[5546] = "test_data_5546.txt";
test_data_files[5547] = "test_data_5547.txt";
test_data_files[5548] = "test_data_5548.txt";
test_data_files[5549] = "test_data_5549.txt";
test_data_files[5550] = "test_data_5550.txt";
test_data_files[5551] = "test_data_5551.txt";
test_data_files[5552] = "test_data_5552.txt";
test_data_files[5553] = "test_data_5553.txt";
test_data_files[5554] = "test_data_5554.txt";
test_data_files[5555] = "test_data_5555.txt";
test_data_files[5556] = "test_data_5556.txt";
test_data_files[5557] = "test_data_5557.txt";
test_data_files[5558] = "test_data_5558.txt";
test_data_files[5559] = "test_data_5559.txt";
test_data_files[5560] = "test_data_5560.txt";
test_data_files[5561] = "test_data_5561.txt";
test_data_files[5562] = "test_data_5562.txt";
test_data_files[5563] = "test_data_5563.txt";
test_data_files[5564] = "test_data_5564.txt";
test_data_files[5565] = "test_data_5565.txt";
test_data_files[5566] = "test_data_5566.txt";
test_data_files[5567] = "test_data_5567.txt";
test_data_files[5568] = "test_data_5568.txt";
test_data_files[5569] = "test_data_5569.txt";
test_data_files[5570] = "test_data_5570.txt";
test_data_files[5571] = "test_data_5571.txt";
test_data_files[5572] = "test_data_5572.txt";
test_data_files[5573] = "test_data_5573.txt";
test_data_files[5574] = "test_data_5574.txt";
test_data_files[5575] = "test_data_5575.txt";
test_data_files[5576] = "test_data_5576.txt";
test_data_files[5577] = "test_data_5577.txt";
test_data_files[5578] = "test_data_5578.txt";
test_data_files[5579] = "test_data_5579.txt";
test_data_files[5580] = "test_data_5580.txt";
test_data_files[5581] = "test_data_5581.txt";
test_data_files[5582] = "test_data_5582.txt";
test_data_files[5583] = "test_data_5583.txt";
test_data_files[5584] = "test_data_5584.txt";
test_data_files[5585] = "test_data_5585.txt";
test_data_files[5586] = "test_data_5586.txt";
test_data_files[5587] = "test_data_5587.txt";
test_data_files[5588] = "test_data_5588.txt";
test_data_files[5589] = "test_data_5589.txt";
test_data_files[5590] = "test_data_5590.txt";
test_data_files[5591] = "test_data_5591.txt";
test_data_files[5592] = "test_data_5592.txt";
test_data_files[5593] = "test_data_5593.txt";
test_data_files[5594] = "test_data_5594.txt";
test_data_files[5595] = "test_data_5595.txt";
test_data_files[5596] = "test_data_5596.txt";
test_data_files[5597] = "test_data_5597.txt";
test_data_files[5598] = "test_data_5598.txt";
test_data_files[5599] = "test_data_5599.txt";
test_data_files[5600] = "test_data_5600.txt";
test_data_files[5601] = "test_data_5601.txt";
test_data_files[5602] = "test_data_5602.txt";
test_data_files[5603] = "test_data_5603.txt";
test_data_files[5604] = "test_data_5604.txt";
test_data_files[5605] = "test_data_5605.txt";
test_data_files[5606] = "test_data_5606.txt";
test_data_files[5607] = "test_data_5607.txt";
test_data_files[5608] = "test_data_5608.txt";
test_data_files[5609] = "test_data_5609.txt";
test_data_files[5610] = "test_data_5610.txt";
test_data_files[5611] = "test_data_5611.txt";
test_data_files[5612] = "test_data_5612.txt";
test_data_files[5613] = "test_data_5613.txt";
test_data_files[5614] = "test_data_5614.txt";
test_data_files[5615] = "test_data_5615.txt";
test_data_files[5616] = "test_data_5616.txt";
test_data_files[5617] = "test_data_5617.txt";
test_data_files[5618] = "test_data_5618.txt";
test_data_files[5619] = "test_data_5619.txt";
test_data_files[5620] = "test_data_5620.txt";
test_data_files[5621] = "test_data_5621.txt";
test_data_files[5622] = "test_data_5622.txt";
test_data_files[5623] = "test_data_5623.txt";
test_data_files[5624] = "test_data_5624.txt";
test_data_files[5625] = "test_data_5625.txt";
test_data_files[5626] = "test_data_5626.txt";
test_data_files[5627] = "test_data_5627.txt";
test_data_files[5628] = "test_data_5628.txt";
test_data_files[5629] = "test_data_5629.txt";
test_data_files[5630] = "test_data_5630.txt";
test_data_files[5631] = "test_data_5631.txt";
test_data_files[5632] = "test_data_5632.txt";
test_data_files[5633] = "test_data_5633.txt";
test_data_files[5634] = "test_data_5634.txt";
test_data_files[5635] = "test_data_5635.txt";
test_data_files[5636] = "test_data_5636.txt";
test_data_files[5637] = "test_data_5637.txt";
test_data_files[5638] = "test_data_5638.txt";
test_data_files[5639] = "test_data_5639.txt";
test_data_files[5640] = "test_data_5640.txt";
test_data_files[5641] = "test_data_5641.txt";
test_data_files[5642] = "test_data_5642.txt";
test_data_files[5643] = "test_data_5643.txt";
test_data_files[5644] = "test_data_5644.txt";
test_data_files[5645] = "test_data_5645.txt";
test_data_files[5646] = "test_data_5646.txt";
test_data_files[5647] = "test_data_5647.txt";
test_data_files[5648] = "test_data_5648.txt";
test_data_files[5649] = "test_data_5649.txt";
test_data_files[5650] = "test_data_5650.txt";
test_data_files[5651] = "test_data_5651.txt";
test_data_files[5652] = "test_data_5652.txt";
test_data_files[5653] = "test_data_5653.txt";
test_data_files[5654] = "test_data_5654.txt";
test_data_files[5655] = "test_data_5655.txt";
test_data_files[5656] = "test_data_5656.txt";
test_data_files[5657] = "test_data_5657.txt";
test_data_files[5658] = "test_data_5658.txt";
test_data_files[5659] = "test_data_5659.txt";
test_data_files[5660] = "test_data_5660.txt";
test_data_files[5661] = "test_data_5661.txt";
test_data_files[5662] = "test_data_5662.txt";
test_data_files[5663] = "test_data_5663.txt";
test_data_files[5664] = "test_data_5664.txt";
test_data_files[5665] = "test_data_5665.txt";
test_data_files[5666] = "test_data_5666.txt";
test_data_files[5667] = "test_data_5667.txt";
test_data_files[5668] = "test_data_5668.txt";
test_data_files[5669] = "test_data_5669.txt";
test_data_files[5670] = "test_data_5670.txt";
test_data_files[5671] = "test_data_5671.txt";
test_data_files[5672] = "test_data_5672.txt";
test_data_files[5673] = "test_data_5673.txt";
test_data_files[5674] = "test_data_5674.txt";
test_data_files[5675] = "test_data_5675.txt";
test_data_files[5676] = "test_data_5676.txt";
test_data_files[5677] = "test_data_5677.txt";
test_data_files[5678] = "test_data_5678.txt";
test_data_files[5679] = "test_data_5679.txt";
test_data_files[5680] = "test_data_5680.txt";
test_data_files[5681] = "test_data_5681.txt";
test_data_files[5682] = "test_data_5682.txt";
test_data_files[5683] = "test_data_5683.txt";
test_data_files[5684] = "test_data_5684.txt";
test_data_files[5685] = "test_data_5685.txt";
test_data_files[5686] = "test_data_5686.txt";
test_data_files[5687] = "test_data_5687.txt";
test_data_files[5688] = "test_data_5688.txt";
test_data_files[5689] = "test_data_5689.txt";
test_data_files[5690] = "test_data_5690.txt";
test_data_files[5691] = "test_data_5691.txt";
test_data_files[5692] = "test_data_5692.txt";
test_data_files[5693] = "test_data_5693.txt";
test_data_files[5694] = "test_data_5694.txt";
test_data_files[5695] = "test_data_5695.txt";
test_data_files[5696] = "test_data_5696.txt";
test_data_files[5697] = "test_data_5697.txt";
test_data_files[5698] = "test_data_5698.txt";
test_data_files[5699] = "test_data_5699.txt";
test_data_files[5700] = "test_data_5700.txt";
test_data_files[5701] = "test_data_5701.txt";
test_data_files[5702] = "test_data_5702.txt";
test_data_files[5703] = "test_data_5703.txt";
test_data_files[5704] = "test_data_5704.txt";
test_data_files[5705] = "test_data_5705.txt";
test_data_files[5706] = "test_data_5706.txt";
test_data_files[5707] = "test_data_5707.txt";
test_data_files[5708] = "test_data_5708.txt";
test_data_files[5709] = "test_data_5709.txt";
test_data_files[5710] = "test_data_5710.txt";
test_data_files[5711] = "test_data_5711.txt";
test_data_files[5712] = "test_data_5712.txt";
test_data_files[5713] = "test_data_5713.txt";
test_data_files[5714] = "test_data_5714.txt";
test_data_files[5715] = "test_data_5715.txt";
test_data_files[5716] = "test_data_5716.txt";
test_data_files[5717] = "test_data_5717.txt";
test_data_files[5718] = "test_data_5718.txt";
test_data_files[5719] = "test_data_5719.txt";
test_data_files[5720] = "test_data_5720.txt";
test_data_files[5721] = "test_data_5721.txt";
test_data_files[5722] = "test_data_5722.txt";
test_data_files[5723] = "test_data_5723.txt";
test_data_files[5724] = "test_data_5724.txt";
test_data_files[5725] = "test_data_5725.txt";
test_data_files[5726] = "test_data_5726.txt";
test_data_files[5727] = "test_data_5727.txt";
test_data_files[5728] = "test_data_5728.txt";
test_data_files[5729] = "test_data_5729.txt";
test_data_files[5730] = "test_data_5730.txt";
test_data_files[5731] = "test_data_5731.txt";
test_data_files[5732] = "test_data_5732.txt";
test_data_files[5733] = "test_data_5733.txt";
test_data_files[5734] = "test_data_5734.txt";
test_data_files[5735] = "test_data_5735.txt";
test_data_files[5736] = "test_data_5736.txt";
test_data_files[5737] = "test_data_5737.txt";
test_data_files[5738] = "test_data_5738.txt";
test_data_files[5739] = "test_data_5739.txt";
test_data_files[5740] = "test_data_5740.txt";
test_data_files[5741] = "test_data_5741.txt";
test_data_files[5742] = "test_data_5742.txt";
test_data_files[5743] = "test_data_5743.txt";
test_data_files[5744] = "test_data_5744.txt";
test_data_files[5745] = "test_data_5745.txt";
test_data_files[5746] = "test_data_5746.txt";
test_data_files[5747] = "test_data_5747.txt";
test_data_files[5748] = "test_data_5748.txt";
test_data_files[5749] = "test_data_5749.txt";
test_data_files[5750] = "test_data_5750.txt";
test_data_files[5751] = "test_data_5751.txt";
test_data_files[5752] = "test_data_5752.txt";
test_data_files[5753] = "test_data_5753.txt";
test_data_files[5754] = "test_data_5754.txt";
test_data_files[5755] = "test_data_5755.txt";
test_data_files[5756] = "test_data_5756.txt";
test_data_files[5757] = "test_data_5757.txt";
test_data_files[5758] = "test_data_5758.txt";
test_data_files[5759] = "test_data_5759.txt";
test_data_files[5760] = "test_data_5760.txt";
test_data_files[5761] = "test_data_5761.txt";
test_data_files[5762] = "test_data_5762.txt";
test_data_files[5763] = "test_data_5763.txt";
test_data_files[5764] = "test_data_5764.txt";
test_data_files[5765] = "test_data_5765.txt";
test_data_files[5766] = "test_data_5766.txt";
test_data_files[5767] = "test_data_5767.txt";
test_data_files[5768] = "test_data_5768.txt";
test_data_files[5769] = "test_data_5769.txt";
test_data_files[5770] = "test_data_5770.txt";
test_data_files[5771] = "test_data_5771.txt";
test_data_files[5772] = "test_data_5772.txt";
test_data_files[5773] = "test_data_5773.txt";
test_data_files[5774] = "test_data_5774.txt";
test_data_files[5775] = "test_data_5775.txt";
test_data_files[5776] = "test_data_5776.txt";
test_data_files[5777] = "test_data_5777.txt";
test_data_files[5778] = "test_data_5778.txt";
test_data_files[5779] = "test_data_5779.txt";
test_data_files[5780] = "test_data_5780.txt";
test_data_files[5781] = "test_data_5781.txt";
test_data_files[5782] = "test_data_5782.txt";
test_data_files[5783] = "test_data_5783.txt";
test_data_files[5784] = "test_data_5784.txt";
test_data_files[5785] = "test_data_5785.txt";
test_data_files[5786] = "test_data_5786.txt";
test_data_files[5787] = "test_data_5787.txt";
test_data_files[5788] = "test_data_5788.txt";
test_data_files[5789] = "test_data_5789.txt";
test_data_files[5790] = "test_data_5790.txt";
test_data_files[5791] = "test_data_5791.txt";
test_data_files[5792] = "test_data_5792.txt";
test_data_files[5793] = "test_data_5793.txt";
test_data_files[5794] = "test_data_5794.txt";
test_data_files[5795] = "test_data_5795.txt";
test_data_files[5796] = "test_data_5796.txt";
test_data_files[5797] = "test_data_5797.txt";
test_data_files[5798] = "test_data_5798.txt";
test_data_files[5799] = "test_data_5799.txt";
test_data_files[5800] = "test_data_5800.txt";
test_data_files[5801] = "test_data_5801.txt";
test_data_files[5802] = "test_data_5802.txt";
test_data_files[5803] = "test_data_5803.txt";
test_data_files[5804] = "test_data_5804.txt";
test_data_files[5805] = "test_data_5805.txt";
test_data_files[5806] = "test_data_5806.txt";
test_data_files[5807] = "test_data_5807.txt";
test_data_files[5808] = "test_data_5808.txt";
test_data_files[5809] = "test_data_5809.txt";
test_data_files[5810] = "test_data_5810.txt";
test_data_files[5811] = "test_data_5811.txt";
test_data_files[5812] = "test_data_5812.txt";
test_data_files[5813] = "test_data_5813.txt";
test_data_files[5814] = "test_data_5814.txt";
test_data_files[5815] = "test_data_5815.txt";
test_data_files[5816] = "test_data_5816.txt";
test_data_files[5817] = "test_data_5817.txt";
test_data_files[5818] = "test_data_5818.txt";
test_data_files[5819] = "test_data_5819.txt";
test_data_files[5820] = "test_data_5820.txt";
test_data_files[5821] = "test_data_5821.txt";
test_data_files[5822] = "test_data_5822.txt";
test_data_files[5823] = "test_data_5823.txt";
test_data_files[5824] = "test_data_5824.txt";
test_data_files[5825] = "test_data_5825.txt";
test_data_files[5826] = "test_data_5826.txt";
test_data_files[5827] = "test_data_5827.txt";
test_data_files[5828] = "test_data_5828.txt";
test_data_files[5829] = "test_data_5829.txt";
test_data_files[5830] = "test_data_5830.txt";
test_data_files[5831] = "test_data_5831.txt";
test_data_files[5832] = "test_data_5832.txt";
test_data_files[5833] = "test_data_5833.txt";
test_data_files[5834] = "test_data_5834.txt";
test_data_files[5835] = "test_data_5835.txt";
test_data_files[5836] = "test_data_5836.txt";
test_data_files[5837] = "test_data_5837.txt";
test_data_files[5838] = "test_data_5838.txt";
test_data_files[5839] = "test_data_5839.txt";
test_data_files[5840] = "test_data_5840.txt";
test_data_files[5841] = "test_data_5841.txt";
test_data_files[5842] = "test_data_5842.txt";
test_data_files[5843] = "test_data_5843.txt";
test_data_files[5844] = "test_data_5844.txt";
test_data_files[5845] = "test_data_5845.txt";
test_data_files[5846] = "test_data_5846.txt";
test_data_files[5847] = "test_data_5847.txt";
test_data_files[5848] = "test_data_5848.txt";
test_data_files[5849] = "test_data_5849.txt";
test_data_files[5850] = "test_data_5850.txt";
test_data_files[5851] = "test_data_5851.txt";
test_data_files[5852] = "test_data_5852.txt";
test_data_files[5853] = "test_data_5853.txt";
test_data_files[5854] = "test_data_5854.txt";
test_data_files[5855] = "test_data_5855.txt";
test_data_files[5856] = "test_data_5856.txt";
test_data_files[5857] = "test_data_5857.txt";
test_data_files[5858] = "test_data_5858.txt";
test_data_files[5859] = "test_data_5859.txt";
test_data_files[5860] = "test_data_5860.txt";
test_data_files[5861] = "test_data_5861.txt";
test_data_files[5862] = "test_data_5862.txt";
test_data_files[5863] = "test_data_5863.txt";
test_data_files[5864] = "test_data_5864.txt";
test_data_files[5865] = "test_data_5865.txt";
test_data_files[5866] = "test_data_5866.txt";
test_data_files[5867] = "test_data_5867.txt";
test_data_files[5868] = "test_data_5868.txt";
test_data_files[5869] = "test_data_5869.txt";
test_data_files[5870] = "test_data_5870.txt";
test_data_files[5871] = "test_data_5871.txt";
test_data_files[5872] = "test_data_5872.txt";
test_data_files[5873] = "test_data_5873.txt";
test_data_files[5874] = "test_data_5874.txt";
test_data_files[5875] = "test_data_5875.txt";
test_data_files[5876] = "test_data_5876.txt";
test_data_files[5877] = "test_data_5877.txt";
test_data_files[5878] = "test_data_5878.txt";
test_data_files[5879] = "test_data_5879.txt";
test_data_files[5880] = "test_data_5880.txt";
test_data_files[5881] = "test_data_5881.txt";
test_data_files[5882] = "test_data_5882.txt";
test_data_files[5883] = "test_data_5883.txt";
test_data_files[5884] = "test_data_5884.txt";
test_data_files[5885] = "test_data_5885.txt";
test_data_files[5886] = "test_data_5886.txt";
test_data_files[5887] = "test_data_5887.txt";
test_data_files[5888] = "test_data_5888.txt";
test_data_files[5889] = "test_data_5889.txt";
test_data_files[5890] = "test_data_5890.txt";
test_data_files[5891] = "test_data_5891.txt";
test_data_files[5892] = "test_data_5892.txt";
test_data_files[5893] = "test_data_5893.txt";
test_data_files[5894] = "test_data_5894.txt";
test_data_files[5895] = "test_data_5895.txt";
test_data_files[5896] = "test_data_5896.txt";
test_data_files[5897] = "test_data_5897.txt";
test_data_files[5898] = "test_data_5898.txt";
test_data_files[5899] = "test_data_5899.txt";
test_data_files[5900] = "test_data_5900.txt";
test_data_files[5901] = "test_data_5901.txt";
test_data_files[5902] = "test_data_5902.txt";
test_data_files[5903] = "test_data_5903.txt";
test_data_files[5904] = "test_data_5904.txt";
test_data_files[5905] = "test_data_5905.txt";
test_data_files[5906] = "test_data_5906.txt";
test_data_files[5907] = "test_data_5907.txt";
test_data_files[5908] = "test_data_5908.txt";
test_data_files[5909] = "test_data_5909.txt";
test_data_files[5910] = "test_data_5910.txt";
test_data_files[5911] = "test_data_5911.txt";
test_data_files[5912] = "test_data_5912.txt";
test_data_files[5913] = "test_data_5913.txt";
test_data_files[5914] = "test_data_5914.txt";
test_data_files[5915] = "test_data_5915.txt";
test_data_files[5916] = "test_data_5916.txt";
test_data_files[5917] = "test_data_5917.txt";
test_data_files[5918] = "test_data_5918.txt";
test_data_files[5919] = "test_data_5919.txt";
test_data_files[5920] = "test_data_5920.txt";
test_data_files[5921] = "test_data_5921.txt";
test_data_files[5922] = "test_data_5922.txt";
test_data_files[5923] = "test_data_5923.txt";
test_data_files[5924] = "test_data_5924.txt";
test_data_files[5925] = "test_data_5925.txt";
test_data_files[5926] = "test_data_5926.txt";
test_data_files[5927] = "test_data_5927.txt";
test_data_files[5928] = "test_data_5928.txt";
test_data_files[5929] = "test_data_5929.txt";
test_data_files[5930] = "test_data_5930.txt";
test_data_files[5931] = "test_data_5931.txt";
test_data_files[5932] = "test_data_5932.txt";
test_data_files[5933] = "test_data_5933.txt";
test_data_files[5934] = "test_data_5934.txt";
test_data_files[5935] = "test_data_5935.txt";
test_data_files[5936] = "test_data_5936.txt";
test_data_files[5937] = "test_data_5937.txt";
test_data_files[5938] = "test_data_5938.txt";
test_data_files[5939] = "test_data_5939.txt";
test_data_files[5940] = "test_data_5940.txt";
test_data_files[5941] = "test_data_5941.txt";
test_data_files[5942] = "test_data_5942.txt";
test_data_files[5943] = "test_data_5943.txt";
test_data_files[5944] = "test_data_5944.txt";
test_data_files[5945] = "test_data_5945.txt";
test_data_files[5946] = "test_data_5946.txt";
test_data_files[5947] = "test_data_5947.txt";
test_data_files[5948] = "test_data_5948.txt";
test_data_files[5949] = "test_data_5949.txt";
test_data_files[5950] = "test_data_5950.txt";
test_data_files[5951] = "test_data_5951.txt";
test_data_files[5952] = "test_data_5952.txt";
test_data_files[5953] = "test_data_5953.txt";
test_data_files[5954] = "test_data_5954.txt";
test_data_files[5955] = "test_data_5955.txt";
test_data_files[5956] = "test_data_5956.txt";
test_data_files[5957] = "test_data_5957.txt";
test_data_files[5958] = "test_data_5958.txt";
test_data_files[5959] = "test_data_5959.txt";
test_data_files[5960] = "test_data_5960.txt";
test_data_files[5961] = "test_data_5961.txt";
test_data_files[5962] = "test_data_5962.txt";
test_data_files[5963] = "test_data_5963.txt";
test_data_files[5964] = "test_data_5964.txt";
test_data_files[5965] = "test_data_5965.txt";
test_data_files[5966] = "test_data_5966.txt";
test_data_files[5967] = "test_data_5967.txt";
test_data_files[5968] = "test_data_5968.txt";
test_data_files[5969] = "test_data_5969.txt";
test_data_files[5970] = "test_data_5970.txt";
test_data_files[5971] = "test_data_5971.txt";
test_data_files[5972] = "test_data_5972.txt";
test_data_files[5973] = "test_data_5973.txt";
test_data_files[5974] = "test_data_5974.txt";
test_data_files[5975] = "test_data_5975.txt";
test_data_files[5976] = "test_data_5976.txt";
test_data_files[5977] = "test_data_5977.txt";
test_data_files[5978] = "test_data_5978.txt";
test_data_files[5979] = "test_data_5979.txt";
test_data_files[5980] = "test_data_5980.txt";
test_data_files[5981] = "test_data_5981.txt";
test_data_files[5982] = "test_data_5982.txt";
test_data_files[5983] = "test_data_5983.txt";
test_data_files[5984] = "test_data_5984.txt";
test_data_files[5985] = "test_data_5985.txt";
test_data_files[5986] = "test_data_5986.txt";
test_data_files[5987] = "test_data_5987.txt";
test_data_files[5988] = "test_data_5988.txt";
test_data_files[5989] = "test_data_5989.txt";
test_data_files[5990] = "test_data_5990.txt";
test_data_files[5991] = "test_data_5991.txt";
test_data_files[5992] = "test_data_5992.txt";
test_data_files[5993] = "test_data_5993.txt";
test_data_files[5994] = "test_data_5994.txt";
test_data_files[5995] = "test_data_5995.txt";
test_data_files[5996] = "test_data_5996.txt";
test_data_files[5997] = "test_data_5997.txt";
test_data_files[5998] = "test_data_5998.txt";
test_data_files[5999] = "test_data_5999.txt";
test_data_files[6000] = "test_data_6000.txt";
test_data_files[6001] = "test_data_6001.txt";
test_data_files[6002] = "test_data_6002.txt";
test_data_files[6003] = "test_data_6003.txt";
test_data_files[6004] = "test_data_6004.txt";
test_data_files[6005] = "test_data_6005.txt";
test_data_files[6006] = "test_data_6006.txt";
test_data_files[6007] = "test_data_6007.txt";
test_data_files[6008] = "test_data_6008.txt";
test_data_files[6009] = "test_data_6009.txt";
test_data_files[6010] = "test_data_6010.txt";
test_data_files[6011] = "test_data_6011.txt";
test_data_files[6012] = "test_data_6012.txt";
test_data_files[6013] = "test_data_6013.txt";
test_data_files[6014] = "test_data_6014.txt";
test_data_files[6015] = "test_data_6015.txt";
test_data_files[6016] = "test_data_6016.txt";
test_data_files[6017] = "test_data_6017.txt";
test_data_files[6018] = "test_data_6018.txt";
test_data_files[6019] = "test_data_6019.txt";
test_data_files[6020] = "test_data_6020.txt";
test_data_files[6021] = "test_data_6021.txt";
test_data_files[6022] = "test_data_6022.txt";
test_data_files[6023] = "test_data_6023.txt";
test_data_files[6024] = "test_data_6024.txt";
test_data_files[6025] = "test_data_6025.txt";
test_data_files[6026] = "test_data_6026.txt";
test_data_files[6027] = "test_data_6027.txt";
test_data_files[6028] = "test_data_6028.txt";
test_data_files[6029] = "test_data_6029.txt";
test_data_files[6030] = "test_data_6030.txt";
test_data_files[6031] = "test_data_6031.txt";
test_data_files[6032] = "test_data_6032.txt";
test_data_files[6033] = "test_data_6033.txt";
test_data_files[6034] = "test_data_6034.txt";
test_data_files[6035] = "test_data_6035.txt";
test_data_files[6036] = "test_data_6036.txt";
test_data_files[6037] = "test_data_6037.txt";
test_data_files[6038] = "test_data_6038.txt";
test_data_files[6039] = "test_data_6039.txt";
test_data_files[6040] = "test_data_6040.txt";
test_data_files[6041] = "test_data_6041.txt";
test_data_files[6042] = "test_data_6042.txt";
test_data_files[6043] = "test_data_6043.txt";
test_data_files[6044] = "test_data_6044.txt";
test_data_files[6045] = "test_data_6045.txt";
test_data_files[6046] = "test_data_6046.txt";
test_data_files[6047] = "test_data_6047.txt";
test_data_files[6048] = "test_data_6048.txt";
test_data_files[6049] = "test_data_6049.txt";
test_data_files[6050] = "test_data_6050.txt";
test_data_files[6051] = "test_data_6051.txt";
test_data_files[6052] = "test_data_6052.txt";
test_data_files[6053] = "test_data_6053.txt";
test_data_files[6054] = "test_data_6054.txt";
test_data_files[6055] = "test_data_6055.txt";
test_data_files[6056] = "test_data_6056.txt";
test_data_files[6057] = "test_data_6057.txt";
test_data_files[6058] = "test_data_6058.txt";
test_data_files[6059] = "test_data_6059.txt";
test_data_files[6060] = "test_data_6060.txt";
test_data_files[6061] = "test_data_6061.txt";
test_data_files[6062] = "test_data_6062.txt";
test_data_files[6063] = "test_data_6063.txt";
test_data_files[6064] = "test_data_6064.txt";
test_data_files[6065] = "test_data_6065.txt";
test_data_files[6066] = "test_data_6066.txt";
test_data_files[6067] = "test_data_6067.txt";
test_data_files[6068] = "test_data_6068.txt";
test_data_files[6069] = "test_data_6069.txt";
test_data_files[6070] = "test_data_6070.txt";
test_data_files[6071] = "test_data_6071.txt";
test_data_files[6072] = "test_data_6072.txt";
test_data_files[6073] = "test_data_6073.txt";
test_data_files[6074] = "test_data_6074.txt";
test_data_files[6075] = "test_data_6075.txt";
test_data_files[6076] = "test_data_6076.txt";
test_data_files[6077] = "test_data_6077.txt";
test_data_files[6078] = "test_data_6078.txt";
test_data_files[6079] = "test_data_6079.txt";
test_data_files[6080] = "test_data_6080.txt";
test_data_files[6081] = "test_data_6081.txt";
test_data_files[6082] = "test_data_6082.txt";
test_data_files[6083] = "test_data_6083.txt";
test_data_files[6084] = "test_data_6084.txt";
test_data_files[6085] = "test_data_6085.txt";
test_data_files[6086] = "test_data_6086.txt";
test_data_files[6087] = "test_data_6087.txt";
test_data_files[6088] = "test_data_6088.txt";
test_data_files[6089] = "test_data_6089.txt";
test_data_files[6090] = "test_data_6090.txt";
test_data_files[6091] = "test_data_6091.txt";
test_data_files[6092] = "test_data_6092.txt";
test_data_files[6093] = "test_data_6093.txt";
test_data_files[6094] = "test_data_6094.txt";
test_data_files[6095] = "test_data_6095.txt";
test_data_files[6096] = "test_data_6096.txt";
test_data_files[6097] = "test_data_6097.txt";
test_data_files[6098] = "test_data_6098.txt";
test_data_files[6099] = "test_data_6099.txt";
test_data_files[6100] = "test_data_6100.txt";
test_data_files[6101] = "test_data_6101.txt";
test_data_files[6102] = "test_data_6102.txt";
test_data_files[6103] = "test_data_6103.txt";
test_data_files[6104] = "test_data_6104.txt";
test_data_files[6105] = "test_data_6105.txt";
test_data_files[6106] = "test_data_6106.txt";
test_data_files[6107] = "test_data_6107.txt";
test_data_files[6108] = "test_data_6108.txt";
test_data_files[6109] = "test_data_6109.txt";
test_data_files[6110] = "test_data_6110.txt";
test_data_files[6111] = "test_data_6111.txt";
test_data_files[6112] = "test_data_6112.txt";
test_data_files[6113] = "test_data_6113.txt";
test_data_files[6114] = "test_data_6114.txt";
test_data_files[6115] = "test_data_6115.txt";
test_data_files[6116] = "test_data_6116.txt";
test_data_files[6117] = "test_data_6117.txt";
test_data_files[6118] = "test_data_6118.txt";
test_data_files[6119] = "test_data_6119.txt";
test_data_files[6120] = "test_data_6120.txt";
test_data_files[6121] = "test_data_6121.txt";
test_data_files[6122] = "test_data_6122.txt";
test_data_files[6123] = "test_data_6123.txt";
test_data_files[6124] = "test_data_6124.txt";
test_data_files[6125] = "test_data_6125.txt";
test_data_files[6126] = "test_data_6126.txt";
test_data_files[6127] = "test_data_6127.txt";
test_data_files[6128] = "test_data_6128.txt";
test_data_files[6129] = "test_data_6129.txt";
test_data_files[6130] = "test_data_6130.txt";
test_data_files[6131] = "test_data_6131.txt";
test_data_files[6132] = "test_data_6132.txt";
test_data_files[6133] = "test_data_6133.txt";
test_data_files[6134] = "test_data_6134.txt";
test_data_files[6135] = "test_data_6135.txt";
test_data_files[6136] = "test_data_6136.txt";
test_data_files[6137] = "test_data_6137.txt";
test_data_files[6138] = "test_data_6138.txt";
test_data_files[6139] = "test_data_6139.txt";
test_data_files[6140] = "test_data_6140.txt";
test_data_files[6141] = "test_data_6141.txt";
test_data_files[6142] = "test_data_6142.txt";
test_data_files[6143] = "test_data_6143.txt";
test_data_files[6144] = "test_data_6144.txt";
test_data_files[6145] = "test_data_6145.txt";
test_data_files[6146] = "test_data_6146.txt";
test_data_files[6147] = "test_data_6147.txt";
test_data_files[6148] = "test_data_6148.txt";
test_data_files[6149] = "test_data_6149.txt";
test_data_files[6150] = "test_data_6150.txt";
test_data_files[6151] = "test_data_6151.txt";
test_data_files[6152] = "test_data_6152.txt";
test_data_files[6153] = "test_data_6153.txt";
test_data_files[6154] = "test_data_6154.txt";
test_data_files[6155] = "test_data_6155.txt";
test_data_files[6156] = "test_data_6156.txt";
test_data_files[6157] = "test_data_6157.txt";
test_data_files[6158] = "test_data_6158.txt";
test_data_files[6159] = "test_data_6159.txt";
test_data_files[6160] = "test_data_6160.txt";
test_data_files[6161] = "test_data_6161.txt";
test_data_files[6162] = "test_data_6162.txt";
test_data_files[6163] = "test_data_6163.txt";
test_data_files[6164] = "test_data_6164.txt";
test_data_files[6165] = "test_data_6165.txt";
test_data_files[6166] = "test_data_6166.txt";
test_data_files[6167] = "test_data_6167.txt";
test_data_files[6168] = "test_data_6168.txt";
test_data_files[6169] = "test_data_6169.txt";
test_data_files[6170] = "test_data_6170.txt";
test_data_files[6171] = "test_data_6171.txt";
test_data_files[6172] = "test_data_6172.txt";
test_data_files[6173] = "test_data_6173.txt";
test_data_files[6174] = "test_data_6174.txt";
test_data_files[6175] = "test_data_6175.txt";
test_data_files[6176] = "test_data_6176.txt";
test_data_files[6177] = "test_data_6177.txt";
test_data_files[6178] = "test_data_6178.txt";
test_data_files[6179] = "test_data_6179.txt";
test_data_files[6180] = "test_data_6180.txt";
test_data_files[6181] = "test_data_6181.txt";
test_data_files[6182] = "test_data_6182.txt";
test_data_files[6183] = "test_data_6183.txt";
test_data_files[6184] = "test_data_6184.txt";
test_data_files[6185] = "test_data_6185.txt";
test_data_files[6186] = "test_data_6186.txt";
test_data_files[6187] = "test_data_6187.txt";
test_data_files[6188] = "test_data_6188.txt";
test_data_files[6189] = "test_data_6189.txt";
test_data_files[6190] = "test_data_6190.txt";
test_data_files[6191] = "test_data_6191.txt";
test_data_files[6192] = "test_data_6192.txt";
test_data_files[6193] = "test_data_6193.txt";
test_data_files[6194] = "test_data_6194.txt";
test_data_files[6195] = "test_data_6195.txt";
test_data_files[6196] = "test_data_6196.txt";
test_data_files[6197] = "test_data_6197.txt";
test_data_files[6198] = "test_data_6198.txt";
test_data_files[6199] = "test_data_6199.txt";
test_data_files[6200] = "test_data_6200.txt";
test_data_files[6201] = "test_data_6201.txt";
test_data_files[6202] = "test_data_6202.txt";
test_data_files[6203] = "test_data_6203.txt";
test_data_files[6204] = "test_data_6204.txt";
test_data_files[6205] = "test_data_6205.txt";
test_data_files[6206] = "test_data_6206.txt";
test_data_files[6207] = "test_data_6207.txt";
test_data_files[6208] = "test_data_6208.txt";
test_data_files[6209] = "test_data_6209.txt";
test_data_files[6210] = "test_data_6210.txt";
test_data_files[6211] = "test_data_6211.txt";
test_data_files[6212] = "test_data_6212.txt";
test_data_files[6213] = "test_data_6213.txt";
test_data_files[6214] = "test_data_6214.txt";
test_data_files[6215] = "test_data_6215.txt";
test_data_files[6216] = "test_data_6216.txt";
test_data_files[6217] = "test_data_6217.txt";
test_data_files[6218] = "test_data_6218.txt";
test_data_files[6219] = "test_data_6219.txt";
test_data_files[6220] = "test_data_6220.txt";
test_data_files[6221] = "test_data_6221.txt";
test_data_files[6222] = "test_data_6222.txt";
test_data_files[6223] = "test_data_6223.txt";
test_data_files[6224] = "test_data_6224.txt";
test_data_files[6225] = "test_data_6225.txt";
test_data_files[6226] = "test_data_6226.txt";
test_data_files[6227] = "test_data_6227.txt";
test_data_files[6228] = "test_data_6228.txt";
test_data_files[6229] = "test_data_6229.txt";
test_data_files[6230] = "test_data_6230.txt";
test_data_files[6231] = "test_data_6231.txt";
test_data_files[6232] = "test_data_6232.txt";
test_data_files[6233] = "test_data_6233.txt";
test_data_files[6234] = "test_data_6234.txt";
test_data_files[6235] = "test_data_6235.txt";
test_data_files[6236] = "test_data_6236.txt";
test_data_files[6237] = "test_data_6237.txt";
test_data_files[6238] = "test_data_6238.txt";
test_data_files[6239] = "test_data_6239.txt";
test_data_files[6240] = "test_data_6240.txt";
test_data_files[6241] = "test_data_6241.txt";
test_data_files[6242] = "test_data_6242.txt";
test_data_files[6243] = "test_data_6243.txt";
test_data_files[6244] = "test_data_6244.txt";
test_data_files[6245] = "test_data_6245.txt";
test_data_files[6246] = "test_data_6246.txt";
test_data_files[6247] = "test_data_6247.txt";
test_data_files[6248] = "test_data_6248.txt";
test_data_files[6249] = "test_data_6249.txt";
test_data_files[6250] = "test_data_6250.txt";
test_data_files[6251] = "test_data_6251.txt";
test_data_files[6252] = "test_data_6252.txt";
test_data_files[6253] = "test_data_6253.txt";
test_data_files[6254] = "test_data_6254.txt";
test_data_files[6255] = "test_data_6255.txt";
test_data_files[6256] = "test_data_6256.txt";
test_data_files[6257] = "test_data_6257.txt";
test_data_files[6258] = "test_data_6258.txt";
test_data_files[6259] = "test_data_6259.txt";
test_data_files[6260] = "test_data_6260.txt";
test_data_files[6261] = "test_data_6261.txt";
test_data_files[6262] = "test_data_6262.txt";
test_data_files[6263] = "test_data_6263.txt";
test_data_files[6264] = "test_data_6264.txt";
test_data_files[6265] = "test_data_6265.txt";
test_data_files[6266] = "test_data_6266.txt";
test_data_files[6267] = "test_data_6267.txt";
test_data_files[6268] = "test_data_6268.txt";
test_data_files[6269] = "test_data_6269.txt";
test_data_files[6270] = "test_data_6270.txt";
test_data_files[6271] = "test_data_6271.txt";
test_data_files[6272] = "test_data_6272.txt";
test_data_files[6273] = "test_data_6273.txt";
test_data_files[6274] = "test_data_6274.txt";
test_data_files[6275] = "test_data_6275.txt";
test_data_files[6276] = "test_data_6276.txt";
test_data_files[6277] = "test_data_6277.txt";
test_data_files[6278] = "test_data_6278.txt";
test_data_files[6279] = "test_data_6279.txt";
test_data_files[6280] = "test_data_6280.txt";
test_data_files[6281] = "test_data_6281.txt";
test_data_files[6282] = "test_data_6282.txt";
test_data_files[6283] = "test_data_6283.txt";
test_data_files[6284] = "test_data_6284.txt";
test_data_files[6285] = "test_data_6285.txt";
test_data_files[6286] = "test_data_6286.txt";
test_data_files[6287] = "test_data_6287.txt";
test_data_files[6288] = "test_data_6288.txt";
test_data_files[6289] = "test_data_6289.txt";
test_data_files[6290] = "test_data_6290.txt";
test_data_files[6291] = "test_data_6291.txt";
test_data_files[6292] = "test_data_6292.txt";
test_data_files[6293] = "test_data_6293.txt";
test_data_files[6294] = "test_data_6294.txt";
test_data_files[6295] = "test_data_6295.txt";
test_data_files[6296] = "test_data_6296.txt";
test_data_files[6297] = "test_data_6297.txt";
test_data_files[6298] = "test_data_6298.txt";
test_data_files[6299] = "test_data_6299.txt";
test_data_files[6300] = "test_data_6300.txt";
test_data_files[6301] = "test_data_6301.txt";
test_data_files[6302] = "test_data_6302.txt";
test_data_files[6303] = "test_data_6303.txt";
test_data_files[6304] = "test_data_6304.txt";
test_data_files[6305] = "test_data_6305.txt";
test_data_files[6306] = "test_data_6306.txt";
test_data_files[6307] = "test_data_6307.txt";
test_data_files[6308] = "test_data_6308.txt";
test_data_files[6309] = "test_data_6309.txt";
test_data_files[6310] = "test_data_6310.txt";
test_data_files[6311] = "test_data_6311.txt";
test_data_files[6312] = "test_data_6312.txt";
test_data_files[6313] = "test_data_6313.txt";
test_data_files[6314] = "test_data_6314.txt";
test_data_files[6315] = "test_data_6315.txt";
test_data_files[6316] = "test_data_6316.txt";
test_data_files[6317] = "test_data_6317.txt";
test_data_files[6318] = "test_data_6318.txt";
test_data_files[6319] = "test_data_6319.txt";
test_data_files[6320] = "test_data_6320.txt";
test_data_files[6321] = "test_data_6321.txt";
test_data_files[6322] = "test_data_6322.txt";
test_data_files[6323] = "test_data_6323.txt";
test_data_files[6324] = "test_data_6324.txt";
test_data_files[6325] = "test_data_6325.txt";
test_data_files[6326] = "test_data_6326.txt";
test_data_files[6327] = "test_data_6327.txt";
test_data_files[6328] = "test_data_6328.txt";
test_data_files[6329] = "test_data_6329.txt";
test_data_files[6330] = "test_data_6330.txt";
test_data_files[6331] = "test_data_6331.txt";
test_data_files[6332] = "test_data_6332.txt";
test_data_files[6333] = "test_data_6333.txt";
test_data_files[6334] = "test_data_6334.txt";
test_data_files[6335] = "test_data_6335.txt";
test_data_files[6336] = "test_data_6336.txt";
test_data_files[6337] = "test_data_6337.txt";
test_data_files[6338] = "test_data_6338.txt";
test_data_files[6339] = "test_data_6339.txt";
test_data_files[6340] = "test_data_6340.txt";
test_data_files[6341] = "test_data_6341.txt";
test_data_files[6342] = "test_data_6342.txt";
test_data_files[6343] = "test_data_6343.txt";
test_data_files[6344] = "test_data_6344.txt";
test_data_files[6345] = "test_data_6345.txt";
test_data_files[6346] = "test_data_6346.txt";
test_data_files[6347] = "test_data_6347.txt";
test_data_files[6348] = "test_data_6348.txt";
test_data_files[6349] = "test_data_6349.txt";
test_data_files[6350] = "test_data_6350.txt";
test_data_files[6351] = "test_data_6351.txt";
test_data_files[6352] = "test_data_6352.txt";
test_data_files[6353] = "test_data_6353.txt";
test_data_files[6354] = "test_data_6354.txt";
test_data_files[6355] = "test_data_6355.txt";
test_data_files[6356] = "test_data_6356.txt";
test_data_files[6357] = "test_data_6357.txt";
test_data_files[6358] = "test_data_6358.txt";
test_data_files[6359] = "test_data_6359.txt";
test_data_files[6360] = "test_data_6360.txt";
test_data_files[6361] = "test_data_6361.txt";
test_data_files[6362] = "test_data_6362.txt";
test_data_files[6363] = "test_data_6363.txt";
test_data_files[6364] = "test_data_6364.txt";
test_data_files[6365] = "test_data_6365.txt";
test_data_files[6366] = "test_data_6366.txt";
test_data_files[6367] = "test_data_6367.txt";
test_data_files[6368] = "test_data_6368.txt";
test_data_files[6369] = "test_data_6369.txt";
test_data_files[6370] = "test_data_6370.txt";
test_data_files[6371] = "test_data_6371.txt";
test_data_files[6372] = "test_data_6372.txt";
test_data_files[6373] = "test_data_6373.txt";
test_data_files[6374] = "test_data_6374.txt";
test_data_files[6375] = "test_data_6375.txt";
test_data_files[6376] = "test_data_6376.txt";
test_data_files[6377] = "test_data_6377.txt";
test_data_files[6378] = "test_data_6378.txt";
test_data_files[6379] = "test_data_6379.txt";
test_data_files[6380] = "test_data_6380.txt";
test_data_files[6381] = "test_data_6381.txt";
test_data_files[6382] = "test_data_6382.txt";
test_data_files[6383] = "test_data_6383.txt";
test_data_files[6384] = "test_data_6384.txt";
test_data_files[6385] = "test_data_6385.txt";
test_data_files[6386] = "test_data_6386.txt";
test_data_files[6387] = "test_data_6387.txt";
test_data_files[6388] = "test_data_6388.txt";
test_data_files[6389] = "test_data_6389.txt";
test_data_files[6390] = "test_data_6390.txt";
test_data_files[6391] = "test_data_6391.txt";
test_data_files[6392] = "test_data_6392.txt";
test_data_files[6393] = "test_data_6393.txt";
test_data_files[6394] = "test_data_6394.txt";
test_data_files[6395] = "test_data_6395.txt";
test_data_files[6396] = "test_data_6396.txt";
test_data_files[6397] = "test_data_6397.txt";
test_data_files[6398] = "test_data_6398.txt";
test_data_files[6399] = "test_data_6399.txt";
test_data_files[6400] = "test_data_6400.txt";
test_data_files[6401] = "test_data_6401.txt";
test_data_files[6402] = "test_data_6402.txt";
test_data_files[6403] = "test_data_6403.txt";
test_data_files[6404] = "test_data_6404.txt";
test_data_files[6405] = "test_data_6405.txt";
test_data_files[6406] = "test_data_6406.txt";
test_data_files[6407] = "test_data_6407.txt";
test_data_files[6408] = "test_data_6408.txt";
test_data_files[6409] = "test_data_6409.txt";
test_data_files[6410] = "test_data_6410.txt";
test_data_files[6411] = "test_data_6411.txt";
test_data_files[6412] = "test_data_6412.txt";
test_data_files[6413] = "test_data_6413.txt";
test_data_files[6414] = "test_data_6414.txt";
test_data_files[6415] = "test_data_6415.txt";
test_data_files[6416] = "test_data_6416.txt";
test_data_files[6417] = "test_data_6417.txt";
test_data_files[6418] = "test_data_6418.txt";
test_data_files[6419] = "test_data_6419.txt";
test_data_files[6420] = "test_data_6420.txt";
test_data_files[6421] = "test_data_6421.txt";
test_data_files[6422] = "test_data_6422.txt";
test_data_files[6423] = "test_data_6423.txt";
test_data_files[6424] = "test_data_6424.txt";
test_data_files[6425] = "test_data_6425.txt";
test_data_files[6426] = "test_data_6426.txt";
test_data_files[6427] = "test_data_6427.txt";
test_data_files[6428] = "test_data_6428.txt";
test_data_files[6429] = "test_data_6429.txt";
test_data_files[6430] = "test_data_6430.txt";
test_data_files[6431] = "test_data_6431.txt";
test_data_files[6432] = "test_data_6432.txt";
test_data_files[6433] = "test_data_6433.txt";
test_data_files[6434] = "test_data_6434.txt";
test_data_files[6435] = "test_data_6435.txt";
test_data_files[6436] = "test_data_6436.txt";
test_data_files[6437] = "test_data_6437.txt";
test_data_files[6438] = "test_data_6438.txt";
test_data_files[6439] = "test_data_6439.txt";
test_data_files[6440] = "test_data_6440.txt";
test_data_files[6441] = "test_data_6441.txt";
test_data_files[6442] = "test_data_6442.txt";
test_data_files[6443] = "test_data_6443.txt";
test_data_files[6444] = "test_data_6444.txt";
test_data_files[6445] = "test_data_6445.txt";
test_data_files[6446] = "test_data_6446.txt";
test_data_files[6447] = "test_data_6447.txt";
test_data_files[6448] = "test_data_6448.txt";
test_data_files[6449] = "test_data_6449.txt";
test_data_files[6450] = "test_data_6450.txt";
test_data_files[6451] = "test_data_6451.txt";
test_data_files[6452] = "test_data_6452.txt";
test_data_files[6453] = "test_data_6453.txt";
test_data_files[6454] = "test_data_6454.txt";
test_data_files[6455] = "test_data_6455.txt";
test_data_files[6456] = "test_data_6456.txt";
test_data_files[6457] = "test_data_6457.txt";
test_data_files[6458] = "test_data_6458.txt";
test_data_files[6459] = "test_data_6459.txt";
test_data_files[6460] = "test_data_6460.txt";
test_data_files[6461] = "test_data_6461.txt";
test_data_files[6462] = "test_data_6462.txt";
test_data_files[6463] = "test_data_6463.txt";
test_data_files[6464] = "test_data_6464.txt";
test_data_files[6465] = "test_data_6465.txt";
test_data_files[6466] = "test_data_6466.txt";
test_data_files[6467] = "test_data_6467.txt";
test_data_files[6468] = "test_data_6468.txt";
test_data_files[6469] = "test_data_6469.txt";
test_data_files[6470] = "test_data_6470.txt";
test_data_files[6471] = "test_data_6471.txt";
test_data_files[6472] = "test_data_6472.txt";
test_data_files[6473] = "test_data_6473.txt";
test_data_files[6474] = "test_data_6474.txt";
test_data_files[6475] = "test_data_6475.txt";
test_data_files[6476] = "test_data_6476.txt";
test_data_files[6477] = "test_data_6477.txt";
test_data_files[6478] = "test_data_6478.txt";
test_data_files[6479] = "test_data_6479.txt";
test_data_files[6480] = "test_data_6480.txt";
test_data_files[6481] = "test_data_6481.txt";
test_data_files[6482] = "test_data_6482.txt";
test_data_files[6483] = "test_data_6483.txt";
test_data_files[6484] = "test_data_6484.txt";
test_data_files[6485] = "test_data_6485.txt";
test_data_files[6486] = "test_data_6486.txt";
test_data_files[6487] = "test_data_6487.txt";
test_data_files[6488] = "test_data_6488.txt";
test_data_files[6489] = "test_data_6489.txt";
test_data_files[6490] = "test_data_6490.txt";
test_data_files[6491] = "test_data_6491.txt";
test_data_files[6492] = "test_data_6492.txt";
test_data_files[6493] = "test_data_6493.txt";
test_data_files[6494] = "test_data_6494.txt";
test_data_files[6495] = "test_data_6495.txt";
test_data_files[6496] = "test_data_6496.txt";
test_data_files[6497] = "test_data_6497.txt";
test_data_files[6498] = "test_data_6498.txt";
test_data_files[6499] = "test_data_6499.txt";
test_data_files[6500] = "test_data_6500.txt";
test_data_files[6501] = "test_data_6501.txt";
test_data_files[6502] = "test_data_6502.txt";
test_data_files[6503] = "test_data_6503.txt";
test_data_files[6504] = "test_data_6504.txt";
test_data_files[6505] = "test_data_6505.txt";
test_data_files[6506] = "test_data_6506.txt";
test_data_files[6507] = "test_data_6507.txt";
test_data_files[6508] = "test_data_6508.txt";
test_data_files[6509] = "test_data_6509.txt";
test_data_files[6510] = "test_data_6510.txt";
test_data_files[6511] = "test_data_6511.txt";
test_data_files[6512] = "test_data_6512.txt";
test_data_files[6513] = "test_data_6513.txt";
test_data_files[6514] = "test_data_6514.txt";
test_data_files[6515] = "test_data_6515.txt";
test_data_files[6516] = "test_data_6516.txt";
test_data_files[6517] = "test_data_6517.txt";
test_data_files[6518] = "test_data_6518.txt";
test_data_files[6519] = "test_data_6519.txt";
test_data_files[6520] = "test_data_6520.txt";
test_data_files[6521] = "test_data_6521.txt";
test_data_files[6522] = "test_data_6522.txt";
test_data_files[6523] = "test_data_6523.txt";
test_data_files[6524] = "test_data_6524.txt";
test_data_files[6525] = "test_data_6525.txt";
test_data_files[6526] = "test_data_6526.txt";
test_data_files[6527] = "test_data_6527.txt";
test_data_files[6528] = "test_data_6528.txt";
test_data_files[6529] = "test_data_6529.txt";
test_data_files[6530] = "test_data_6530.txt";
test_data_files[6531] = "test_data_6531.txt";
test_data_files[6532] = "test_data_6532.txt";
test_data_files[6533] = "test_data_6533.txt";
test_data_files[6534] = "test_data_6534.txt";
test_data_files[6535] = "test_data_6535.txt";
test_data_files[6536] = "test_data_6536.txt";
test_data_files[6537] = "test_data_6537.txt";
test_data_files[6538] = "test_data_6538.txt";
test_data_files[6539] = "test_data_6539.txt";
test_data_files[6540] = "test_data_6540.txt";
test_data_files[6541] = "test_data_6541.txt";
test_data_files[6542] = "test_data_6542.txt";
test_data_files[6543] = "test_data_6543.txt";
test_data_files[6544] = "test_data_6544.txt";
test_data_files[6545] = "test_data_6545.txt";
test_data_files[6546] = "test_data_6546.txt";
test_data_files[6547] = "test_data_6547.txt";
test_data_files[6548] = "test_data_6548.txt";
test_data_files[6549] = "test_data_6549.txt";
test_data_files[6550] = "test_data_6550.txt";
test_data_files[6551] = "test_data_6551.txt";
test_data_files[6552] = "test_data_6552.txt";
test_data_files[6553] = "test_data_6553.txt";
test_data_files[6554] = "test_data_6554.txt";
test_data_files[6555] = "test_data_6555.txt";
test_data_files[6556] = "test_data_6556.txt";
test_data_files[6557] = "test_data_6557.txt";
test_data_files[6558] = "test_data_6558.txt";
test_data_files[6559] = "test_data_6559.txt";
test_data_files[6560] = "test_data_6560.txt";
test_data_files[6561] = "test_data_6561.txt";
test_data_files[6562] = "test_data_6562.txt";
test_data_files[6563] = "test_data_6563.txt";
test_data_files[6564] = "test_data_6564.txt";
test_data_files[6565] = "test_data_6565.txt";
test_data_files[6566] = "test_data_6566.txt";
test_data_files[6567] = "test_data_6567.txt";
test_data_files[6568] = "test_data_6568.txt";
test_data_files[6569] = "test_data_6569.txt";
test_data_files[6570] = "test_data_6570.txt";
test_data_files[6571] = "test_data_6571.txt";
test_data_files[6572] = "test_data_6572.txt";
test_data_files[6573] = "test_data_6573.txt";
test_data_files[6574] = "test_data_6574.txt";
test_data_files[6575] = "test_data_6575.txt";
test_data_files[6576] = "test_data_6576.txt";
test_data_files[6577] = "test_data_6577.txt";
test_data_files[6578] = "test_data_6578.txt";
test_data_files[6579] = "test_data_6579.txt";
test_data_files[6580] = "test_data_6580.txt";
test_data_files[6581] = "test_data_6581.txt";
test_data_files[6582] = "test_data_6582.txt";
test_data_files[6583] = "test_data_6583.txt";
test_data_files[6584] = "test_data_6584.txt";
test_data_files[6585] = "test_data_6585.txt";
test_data_files[6586] = "test_data_6586.txt";
test_data_files[6587] = "test_data_6587.txt";
test_data_files[6588] = "test_data_6588.txt";
test_data_files[6589] = "test_data_6589.txt";
test_data_files[6590] = "test_data_6590.txt";
test_data_files[6591] = "test_data_6591.txt";
test_data_files[6592] = "test_data_6592.txt";
test_data_files[6593] = "test_data_6593.txt";
test_data_files[6594] = "test_data_6594.txt";
test_data_files[6595] = "test_data_6595.txt";
test_data_files[6596] = "test_data_6596.txt";
test_data_files[6597] = "test_data_6597.txt";
test_data_files[6598] = "test_data_6598.txt";
test_data_files[6599] = "test_data_6599.txt";
test_data_files[6600] = "test_data_6600.txt";
test_data_files[6601] = "test_data_6601.txt";
test_data_files[6602] = "test_data_6602.txt";
test_data_files[6603] = "test_data_6603.txt";
test_data_files[6604] = "test_data_6604.txt";
test_data_files[6605] = "test_data_6605.txt";
test_data_files[6606] = "test_data_6606.txt";
test_data_files[6607] = "test_data_6607.txt";
test_data_files[6608] = "test_data_6608.txt";
test_data_files[6609] = "test_data_6609.txt";
test_data_files[6610] = "test_data_6610.txt";
test_data_files[6611] = "test_data_6611.txt";
test_data_files[6612] = "test_data_6612.txt";
test_data_files[6613] = "test_data_6613.txt";
test_data_files[6614] = "test_data_6614.txt";
test_data_files[6615] = "test_data_6615.txt";
test_data_files[6616] = "test_data_6616.txt";
test_data_files[6617] = "test_data_6617.txt";
test_data_files[6618] = "test_data_6618.txt";
test_data_files[6619] = "test_data_6619.txt";
test_data_files[6620] = "test_data_6620.txt";
test_data_files[6621] = "test_data_6621.txt";
test_data_files[6622] = "test_data_6622.txt";
test_data_files[6623] = "test_data_6623.txt";
test_data_files[6624] = "test_data_6624.txt";
test_data_files[6625] = "test_data_6625.txt";
test_data_files[6626] = "test_data_6626.txt";
test_data_files[6627] = "test_data_6627.txt";
test_data_files[6628] = "test_data_6628.txt";
test_data_files[6629] = "test_data_6629.txt";
test_data_files[6630] = "test_data_6630.txt";
test_data_files[6631] = "test_data_6631.txt";
test_data_files[6632] = "test_data_6632.txt";
test_data_files[6633] = "test_data_6633.txt";
test_data_files[6634] = "test_data_6634.txt";
test_data_files[6635] = "test_data_6635.txt";
test_data_files[6636] = "test_data_6636.txt";
test_data_files[6637] = "test_data_6637.txt";
test_data_files[6638] = "test_data_6638.txt";
test_data_files[6639] = "test_data_6639.txt";
test_data_files[6640] = "test_data_6640.txt";
test_data_files[6641] = "test_data_6641.txt";
test_data_files[6642] = "test_data_6642.txt";
test_data_files[6643] = "test_data_6643.txt";
test_data_files[6644] = "test_data_6644.txt";
test_data_files[6645] = "test_data_6645.txt";
test_data_files[6646] = "test_data_6646.txt";
test_data_files[6647] = "test_data_6647.txt";
test_data_files[6648] = "test_data_6648.txt";
test_data_files[6649] = "test_data_6649.txt";
test_data_files[6650] = "test_data_6650.txt";
test_data_files[6651] = "test_data_6651.txt";
test_data_files[6652] = "test_data_6652.txt";
test_data_files[6653] = "test_data_6653.txt";
test_data_files[6654] = "test_data_6654.txt";
test_data_files[6655] = "test_data_6655.txt";
test_data_files[6656] = "test_data_6656.txt";
test_data_files[6657] = "test_data_6657.txt";
test_data_files[6658] = "test_data_6658.txt";
test_data_files[6659] = "test_data_6659.txt";
test_data_files[6660] = "test_data_6660.txt";
test_data_files[6661] = "test_data_6661.txt";
test_data_files[6662] = "test_data_6662.txt";
test_data_files[6663] = "test_data_6663.txt";
test_data_files[6664] = "test_data_6664.txt";
test_data_files[6665] = "test_data_6665.txt";
test_data_files[6666] = "test_data_6666.txt";
test_data_files[6667] = "test_data_6667.txt";
test_data_files[6668] = "test_data_6668.txt";
test_data_files[6669] = "test_data_6669.txt";
test_data_files[6670] = "test_data_6670.txt";
test_data_files[6671] = "test_data_6671.txt";
test_data_files[6672] = "test_data_6672.txt";
test_data_files[6673] = "test_data_6673.txt";
test_data_files[6674] = "test_data_6674.txt";
test_data_files[6675] = "test_data_6675.txt";
test_data_files[6676] = "test_data_6676.txt";
test_data_files[6677] = "test_data_6677.txt";
test_data_files[6678] = "test_data_6678.txt";
test_data_files[6679] = "test_data_6679.txt";
test_data_files[6680] = "test_data_6680.txt";
test_data_files[6681] = "test_data_6681.txt";
test_data_files[6682] = "test_data_6682.txt";
test_data_files[6683] = "test_data_6683.txt";
test_data_files[6684] = "test_data_6684.txt";
test_data_files[6685] = "test_data_6685.txt";
test_data_files[6686] = "test_data_6686.txt";
test_data_files[6687] = "test_data_6687.txt";
test_data_files[6688] = "test_data_6688.txt";
test_data_files[6689] = "test_data_6689.txt";
test_data_files[6690] = "test_data_6690.txt";
test_data_files[6691] = "test_data_6691.txt";
test_data_files[6692] = "test_data_6692.txt";
test_data_files[6693] = "test_data_6693.txt";
test_data_files[6694] = "test_data_6694.txt";
test_data_files[6695] = "test_data_6695.txt";
test_data_files[6696] = "test_data_6696.txt";
test_data_files[6697] = "test_data_6697.txt";
test_data_files[6698] = "test_data_6698.txt";
test_data_files[6699] = "test_data_6699.txt";
test_data_files[6700] = "test_data_6700.txt";
test_data_files[6701] = "test_data_6701.txt";
test_data_files[6702] = "test_data_6702.txt";
test_data_files[6703] = "test_data_6703.txt";
test_data_files[6704] = "test_data_6704.txt";
test_data_files[6705] = "test_data_6705.txt";
test_data_files[6706] = "test_data_6706.txt";
test_data_files[6707] = "test_data_6707.txt";
test_data_files[6708] = "test_data_6708.txt";
test_data_files[6709] = "test_data_6709.txt";
test_data_files[6710] = "test_data_6710.txt";
test_data_files[6711] = "test_data_6711.txt";
test_data_files[6712] = "test_data_6712.txt";
test_data_files[6713] = "test_data_6713.txt";
test_data_files[6714] = "test_data_6714.txt";
test_data_files[6715] = "test_data_6715.txt";
test_data_files[6716] = "test_data_6716.txt";
test_data_files[6717] = "test_data_6717.txt";
test_data_files[6718] = "test_data_6718.txt";
test_data_files[6719] = "test_data_6719.txt";
test_data_files[6720] = "test_data_6720.txt";
test_data_files[6721] = "test_data_6721.txt";
test_data_files[6722] = "test_data_6722.txt";
test_data_files[6723] = "test_data_6723.txt";
test_data_files[6724] = "test_data_6724.txt";
test_data_files[6725] = "test_data_6725.txt";
test_data_files[6726] = "test_data_6726.txt";
test_data_files[6727] = "test_data_6727.txt";
test_data_files[6728] = "test_data_6728.txt";
test_data_files[6729] = "test_data_6729.txt";
test_data_files[6730] = "test_data_6730.txt";
test_data_files[6731] = "test_data_6731.txt";
test_data_files[6732] = "test_data_6732.txt";
test_data_files[6733] = "test_data_6733.txt";
test_data_files[6734] = "test_data_6734.txt";
test_data_files[6735] = "test_data_6735.txt";
test_data_files[6736] = "test_data_6736.txt";
test_data_files[6737] = "test_data_6737.txt";
test_data_files[6738] = "test_data_6738.txt";
test_data_files[6739] = "test_data_6739.txt";
test_data_files[6740] = "test_data_6740.txt";
test_data_files[6741] = "test_data_6741.txt";
test_data_files[6742] = "test_data_6742.txt";
test_data_files[6743] = "test_data_6743.txt";
test_data_files[6744] = "test_data_6744.txt";
test_data_files[6745] = "test_data_6745.txt";
test_data_files[6746] = "test_data_6746.txt";
test_data_files[6747] = "test_data_6747.txt";
test_data_files[6748] = "test_data_6748.txt";
test_data_files[6749] = "test_data_6749.txt";
test_data_files[6750] = "test_data_6750.txt";
test_data_files[6751] = "test_data_6751.txt";
test_data_files[6752] = "test_data_6752.txt";
test_data_files[6753] = "test_data_6753.txt";
test_data_files[6754] = "test_data_6754.txt";
test_data_files[6755] = "test_data_6755.txt";
test_data_files[6756] = "test_data_6756.txt";
test_data_files[6757] = "test_data_6757.txt";
test_data_files[6758] = "test_data_6758.txt";
test_data_files[6759] = "test_data_6759.txt";
test_data_files[6760] = "test_data_6760.txt";
test_data_files[6761] = "test_data_6761.txt";
test_data_files[6762] = "test_data_6762.txt";
test_data_files[6763] = "test_data_6763.txt";
test_data_files[6764] = "test_data_6764.txt";
test_data_files[6765] = "test_data_6765.txt";
test_data_files[6766] = "test_data_6766.txt";
test_data_files[6767] = "test_data_6767.txt";
test_data_files[6768] = "test_data_6768.txt";
test_data_files[6769] = "test_data_6769.txt";
test_data_files[6770] = "test_data_6770.txt";
test_data_files[6771] = "test_data_6771.txt";
test_data_files[6772] = "test_data_6772.txt";
test_data_files[6773] = "test_data_6773.txt";
test_data_files[6774] = "test_data_6774.txt";
test_data_files[6775] = "test_data_6775.txt";
test_data_files[6776] = "test_data_6776.txt";
test_data_files[6777] = "test_data_6777.txt";
test_data_files[6778] = "test_data_6778.txt";
test_data_files[6779] = "test_data_6779.txt";
test_data_files[6780] = "test_data_6780.txt";
test_data_files[6781] = "test_data_6781.txt";
test_data_files[6782] = "test_data_6782.txt";
test_data_files[6783] = "test_data_6783.txt";
test_data_files[6784] = "test_data_6784.txt";
test_data_files[6785] = "test_data_6785.txt";
test_data_files[6786] = "test_data_6786.txt";
test_data_files[6787] = "test_data_6787.txt";
test_data_files[6788] = "test_data_6788.txt";
test_data_files[6789] = "test_data_6789.txt";
test_data_files[6790] = "test_data_6790.txt";
test_data_files[6791] = "test_data_6791.txt";
test_data_files[6792] = "test_data_6792.txt";
test_data_files[6793] = "test_data_6793.txt";
test_data_files[6794] = "test_data_6794.txt";
test_data_files[6795] = "test_data_6795.txt";
test_data_files[6796] = "test_data_6796.txt";
test_data_files[6797] = "test_data_6797.txt";
test_data_files[6798] = "test_data_6798.txt";
test_data_files[6799] = "test_data_6799.txt";
test_data_files[6800] = "test_data_6800.txt";
test_data_files[6801] = "test_data_6801.txt";
test_data_files[6802] = "test_data_6802.txt";
test_data_files[6803] = "test_data_6803.txt";
test_data_files[6804] = "test_data_6804.txt";
test_data_files[6805] = "test_data_6805.txt";
test_data_files[6806] = "test_data_6806.txt";
test_data_files[6807] = "test_data_6807.txt";
test_data_files[6808] = "test_data_6808.txt";
test_data_files[6809] = "test_data_6809.txt";
test_data_files[6810] = "test_data_6810.txt";
test_data_files[6811] = "test_data_6811.txt";
test_data_files[6812] = "test_data_6812.txt";
test_data_files[6813] = "test_data_6813.txt";
test_data_files[6814] = "test_data_6814.txt";
test_data_files[6815] = "test_data_6815.txt";
test_data_files[6816] = "test_data_6816.txt";
test_data_files[6817] = "test_data_6817.txt";
test_data_files[6818] = "test_data_6818.txt";
test_data_files[6819] = "test_data_6819.txt";
test_data_files[6820] = "test_data_6820.txt";
test_data_files[6821] = "test_data_6821.txt";
test_data_files[6822] = "test_data_6822.txt";
test_data_files[6823] = "test_data_6823.txt";
test_data_files[6824] = "test_data_6824.txt";
test_data_files[6825] = "test_data_6825.txt";
test_data_files[6826] = "test_data_6826.txt";
test_data_files[6827] = "test_data_6827.txt";
test_data_files[6828] = "test_data_6828.txt";
test_data_files[6829] = "test_data_6829.txt";
test_data_files[6830] = "test_data_6830.txt";
test_data_files[6831] = "test_data_6831.txt";
test_data_files[6832] = "test_data_6832.txt";
test_data_files[6833] = "test_data_6833.txt";
test_data_files[6834] = "test_data_6834.txt";
test_data_files[6835] = "test_data_6835.txt";
test_data_files[6836] = "test_data_6836.txt";
test_data_files[6837] = "test_data_6837.txt";
test_data_files[6838] = "test_data_6838.txt";
test_data_files[6839] = "test_data_6839.txt";
test_data_files[6840] = "test_data_6840.txt";
test_data_files[6841] = "test_data_6841.txt";
test_data_files[6842] = "test_data_6842.txt";
test_data_files[6843] = "test_data_6843.txt";
test_data_files[6844] = "test_data_6844.txt";
test_data_files[6845] = "test_data_6845.txt";
test_data_files[6846] = "test_data_6846.txt";
test_data_files[6847] = "test_data_6847.txt";
test_data_files[6848] = "test_data_6848.txt";
test_data_files[6849] = "test_data_6849.txt";
test_data_files[6850] = "test_data_6850.txt";
test_data_files[6851] = "test_data_6851.txt";
test_data_files[6852] = "test_data_6852.txt";
test_data_files[6853] = "test_data_6853.txt";
test_data_files[6854] = "test_data_6854.txt";
test_data_files[6855] = "test_data_6855.txt";
test_data_files[6856] = "test_data_6856.txt";
test_data_files[6857] = "test_data_6857.txt";
test_data_files[6858] = "test_data_6858.txt";
test_data_files[6859] = "test_data_6859.txt";
test_data_files[6860] = "test_data_6860.txt";
test_data_files[6861] = "test_data_6861.txt";
test_data_files[6862] = "test_data_6862.txt";
test_data_files[6863] = "test_data_6863.txt";
test_data_files[6864] = "test_data_6864.txt";
test_data_files[6865] = "test_data_6865.txt";
test_data_files[6866] = "test_data_6866.txt";
test_data_files[6867] = "test_data_6867.txt";
test_data_files[6868] = "test_data_6868.txt";
test_data_files[6869] = "test_data_6869.txt";
test_data_files[6870] = "test_data_6870.txt";
test_data_files[6871] = "test_data_6871.txt";
test_data_files[6872] = "test_data_6872.txt";
test_data_files[6873] = "test_data_6873.txt";
test_data_files[6874] = "test_data_6874.txt";
test_data_files[6875] = "test_data_6875.txt";
test_data_files[6876] = "test_data_6876.txt";
test_data_files[6877] = "test_data_6877.txt";
test_data_files[6878] = "test_data_6878.txt";
test_data_files[6879] = "test_data_6879.txt";
test_data_files[6880] = "test_data_6880.txt";
test_data_files[6881] = "test_data_6881.txt";
test_data_files[6882] = "test_data_6882.txt";
test_data_files[6883] = "test_data_6883.txt";
test_data_files[6884] = "test_data_6884.txt";
test_data_files[6885] = "test_data_6885.txt";
test_data_files[6886] = "test_data_6886.txt";
test_data_files[6887] = "test_data_6887.txt";
test_data_files[6888] = "test_data_6888.txt";
test_data_files[6889] = "test_data_6889.txt";
test_data_files[6890] = "test_data_6890.txt";
test_data_files[6891] = "test_data_6891.txt";
test_data_files[6892] = "test_data_6892.txt";
test_data_files[6893] = "test_data_6893.txt";
test_data_files[6894] = "test_data_6894.txt";
test_data_files[6895] = "test_data_6895.txt";
test_data_files[6896] = "test_data_6896.txt";
test_data_files[6897] = "test_data_6897.txt";
test_data_files[6898] = "test_data_6898.txt";
test_data_files[6899] = "test_data_6899.txt";
test_data_files[6900] = "test_data_6900.txt";
test_data_files[6901] = "test_data_6901.txt";
test_data_files[6902] = "test_data_6902.txt";
test_data_files[6903] = "test_data_6903.txt";
test_data_files[6904] = "test_data_6904.txt";
test_data_files[6905] = "test_data_6905.txt";
test_data_files[6906] = "test_data_6906.txt";
test_data_files[6907] = "test_data_6907.txt";
test_data_files[6908] = "test_data_6908.txt";
test_data_files[6909] = "test_data_6909.txt";
test_data_files[6910] = "test_data_6910.txt";
test_data_files[6911] = "test_data_6911.txt";
test_data_files[6912] = "test_data_6912.txt";
test_data_files[6913] = "test_data_6913.txt";
test_data_files[6914] = "test_data_6914.txt";
test_data_files[6915] = "test_data_6915.txt";
test_data_files[6916] = "test_data_6916.txt";
test_data_files[6917] = "test_data_6917.txt";
test_data_files[6918] = "test_data_6918.txt";
test_data_files[6919] = "test_data_6919.txt";
test_data_files[6920] = "test_data_6920.txt";
test_data_files[6921] = "test_data_6921.txt";
test_data_files[6922] = "test_data_6922.txt";
test_data_files[6923] = "test_data_6923.txt";
test_data_files[6924] = "test_data_6924.txt";
test_data_files[6925] = "test_data_6925.txt";
test_data_files[6926] = "test_data_6926.txt";
test_data_files[6927] = "test_data_6927.txt";
test_data_files[6928] = "test_data_6928.txt";
test_data_files[6929] = "test_data_6929.txt";
test_data_files[6930] = "test_data_6930.txt";
test_data_files[6931] = "test_data_6931.txt";
test_data_files[6932] = "test_data_6932.txt";
test_data_files[6933] = "test_data_6933.txt";
test_data_files[6934] = "test_data_6934.txt";
test_data_files[6935] = "test_data_6935.txt";
test_data_files[6936] = "test_data_6936.txt";
test_data_files[6937] = "test_data_6937.txt";
test_data_files[6938] = "test_data_6938.txt";
test_data_files[6939] = "test_data_6939.txt";
test_data_files[6940] = "test_data_6940.txt";
test_data_files[6941] = "test_data_6941.txt";
test_data_files[6942] = "test_data_6942.txt";
test_data_files[6943] = "test_data_6943.txt";
test_data_files[6944] = "test_data_6944.txt";
test_data_files[6945] = "test_data_6945.txt";
test_data_files[6946] = "test_data_6946.txt";
test_data_files[6947] = "test_data_6947.txt";
test_data_files[6948] = "test_data_6948.txt";
test_data_files[6949] = "test_data_6949.txt";
test_data_files[6950] = "test_data_6950.txt";
test_data_files[6951] = "test_data_6951.txt";
test_data_files[6952] = "test_data_6952.txt";
test_data_files[6953] = "test_data_6953.txt";
test_data_files[6954] = "test_data_6954.txt";
test_data_files[6955] = "test_data_6955.txt";
test_data_files[6956] = "test_data_6956.txt";
test_data_files[6957] = "test_data_6957.txt";
test_data_files[6958] = "test_data_6958.txt";
test_data_files[6959] = "test_data_6959.txt";
test_data_files[6960] = "test_data_6960.txt";
test_data_files[6961] = "test_data_6961.txt";
test_data_files[6962] = "test_data_6962.txt";
test_data_files[6963] = "test_data_6963.txt";
test_data_files[6964] = "test_data_6964.txt";
test_data_files[6965] = "test_data_6965.txt";
test_data_files[6966] = "test_data_6966.txt";
test_data_files[6967] = "test_data_6967.txt";
test_data_files[6968] = "test_data_6968.txt";
test_data_files[6969] = "test_data_6969.txt";
test_data_files[6970] = "test_data_6970.txt";
test_data_files[6971] = "test_data_6971.txt";
test_data_files[6972] = "test_data_6972.txt";
test_data_files[6973] = "test_data_6973.txt";
test_data_files[6974] = "test_data_6974.txt";
test_data_files[6975] = "test_data_6975.txt";
test_data_files[6976] = "test_data_6976.txt";
test_data_files[6977] = "test_data_6977.txt";
test_data_files[6978] = "test_data_6978.txt";
test_data_files[6979] = "test_data_6979.txt";
test_data_files[6980] = "test_data_6980.txt";
test_data_files[6981] = "test_data_6981.txt";
test_data_files[6982] = "test_data_6982.txt";
test_data_files[6983] = "test_data_6983.txt";
test_data_files[6984] = "test_data_6984.txt";
test_data_files[6985] = "test_data_6985.txt";
test_data_files[6986] = "test_data_6986.txt";
test_data_files[6987] = "test_data_6987.txt";
test_data_files[6988] = "test_data_6988.txt";
test_data_files[6989] = "test_data_6989.txt";
test_data_files[6990] = "test_data_6990.txt";
test_data_files[6991] = "test_data_6991.txt";
test_data_files[6992] = "test_data_6992.txt";
test_data_files[6993] = "test_data_6993.txt";
test_data_files[6994] = "test_data_6994.txt";
test_data_files[6995] = "test_data_6995.txt";
test_data_files[6996] = "test_data_6996.txt";
test_data_files[6997] = "test_data_6997.txt";
test_data_files[6998] = "test_data_6998.txt";
test_data_files[6999] = "test_data_6999.txt";
test_data_files[7000] = "test_data_7000.txt";
test_data_files[7001] = "test_data_7001.txt";
test_data_files[7002] = "test_data_7002.txt";
test_data_files[7003] = "test_data_7003.txt";
test_data_files[7004] = "test_data_7004.txt";
test_data_files[7005] = "test_data_7005.txt";
test_data_files[7006] = "test_data_7006.txt";
test_data_files[7007] = "test_data_7007.txt";
test_data_files[7008] = "test_data_7008.txt";
test_data_files[7009] = "test_data_7009.txt";
test_data_files[7010] = "test_data_7010.txt";
test_data_files[7011] = "test_data_7011.txt";
test_data_files[7012] = "test_data_7012.txt";
test_data_files[7013] = "test_data_7013.txt";
test_data_files[7014] = "test_data_7014.txt";
test_data_files[7015] = "test_data_7015.txt";
test_data_files[7016] = "test_data_7016.txt";
test_data_files[7017] = "test_data_7017.txt";
test_data_files[7018] = "test_data_7018.txt";
test_data_files[7019] = "test_data_7019.txt";
test_data_files[7020] = "test_data_7020.txt";
test_data_files[7021] = "test_data_7021.txt";
test_data_files[7022] = "test_data_7022.txt";
test_data_files[7023] = "test_data_7023.txt";
test_data_files[7024] = "test_data_7024.txt";
test_data_files[7025] = "test_data_7025.txt";
test_data_files[7026] = "test_data_7026.txt";
test_data_files[7027] = "test_data_7027.txt";
test_data_files[7028] = "test_data_7028.txt";
test_data_files[7029] = "test_data_7029.txt";
test_data_files[7030] = "test_data_7030.txt";
test_data_files[7031] = "test_data_7031.txt";
test_data_files[7032] = "test_data_7032.txt";
test_data_files[7033] = "test_data_7033.txt";
test_data_files[7034] = "test_data_7034.txt";
test_data_files[7035] = "test_data_7035.txt";
test_data_files[7036] = "test_data_7036.txt";
test_data_files[7037] = "test_data_7037.txt";
test_data_files[7038] = "test_data_7038.txt";
test_data_files[7039] = "test_data_7039.txt";
test_data_files[7040] = "test_data_7040.txt";
test_data_files[7041] = "test_data_7041.txt";
test_data_files[7042] = "test_data_7042.txt";
test_data_files[7043] = "test_data_7043.txt";
test_data_files[7044] = "test_data_7044.txt";
test_data_files[7045] = "test_data_7045.txt";
test_data_files[7046] = "test_data_7046.txt";
test_data_files[7047] = "test_data_7047.txt";
test_data_files[7048] = "test_data_7048.txt";
test_data_files[7049] = "test_data_7049.txt";
test_data_files[7050] = "test_data_7050.txt";
test_data_files[7051] = "test_data_7051.txt";
test_data_files[7052] = "test_data_7052.txt";
test_data_files[7053] = "test_data_7053.txt";
test_data_files[7054] = "test_data_7054.txt";
test_data_files[7055] = "test_data_7055.txt";
test_data_files[7056] = "test_data_7056.txt";
test_data_files[7057] = "test_data_7057.txt";
test_data_files[7058] = "test_data_7058.txt";
test_data_files[7059] = "test_data_7059.txt";
test_data_files[7060] = "test_data_7060.txt";
test_data_files[7061] = "test_data_7061.txt";
test_data_files[7062] = "test_data_7062.txt";
test_data_files[7063] = "test_data_7063.txt";
test_data_files[7064] = "test_data_7064.txt";
test_data_files[7065] = "test_data_7065.txt";
test_data_files[7066] = "test_data_7066.txt";
test_data_files[7067] = "test_data_7067.txt";
test_data_files[7068] = "test_data_7068.txt";
test_data_files[7069] = "test_data_7069.txt";
test_data_files[7070] = "test_data_7070.txt";
test_data_files[7071] = "test_data_7071.txt";
test_data_files[7072] = "test_data_7072.txt";
test_data_files[7073] = "test_data_7073.txt";
test_data_files[7074] = "test_data_7074.txt";
test_data_files[7075] = "test_data_7075.txt";
test_data_files[7076] = "test_data_7076.txt";
test_data_files[7077] = "test_data_7077.txt";
test_data_files[7078] = "test_data_7078.txt";
test_data_files[7079] = "test_data_7079.txt";
test_data_files[7080] = "test_data_7080.txt";
test_data_files[7081] = "test_data_7081.txt";
test_data_files[7082] = "test_data_7082.txt";
test_data_files[7083] = "test_data_7083.txt";
test_data_files[7084] = "test_data_7084.txt";
test_data_files[7085] = "test_data_7085.txt";
test_data_files[7086] = "test_data_7086.txt";
test_data_files[7087] = "test_data_7087.txt";
test_data_files[7088] = "test_data_7088.txt";
test_data_files[7089] = "test_data_7089.txt";
test_data_files[7090] = "test_data_7090.txt";
test_data_files[7091] = "test_data_7091.txt";
test_data_files[7092] = "test_data_7092.txt";
test_data_files[7093] = "test_data_7093.txt";
test_data_files[7094] = "test_data_7094.txt";
test_data_files[7095] = "test_data_7095.txt";
test_data_files[7096] = "test_data_7096.txt";
test_data_files[7097] = "test_data_7097.txt";
test_data_files[7098] = "test_data_7098.txt";
test_data_files[7099] = "test_data_7099.txt";
test_data_files[7100] = "test_data_7100.txt";
test_data_files[7101] = "test_data_7101.txt";
test_data_files[7102] = "test_data_7102.txt";
test_data_files[7103] = "test_data_7103.txt";
test_data_files[7104] = "test_data_7104.txt";
test_data_files[7105] = "test_data_7105.txt";
test_data_files[7106] = "test_data_7106.txt";
test_data_files[7107] = "test_data_7107.txt";
test_data_files[7108] = "test_data_7108.txt";
test_data_files[7109] = "test_data_7109.txt";
test_data_files[7110] = "test_data_7110.txt";
test_data_files[7111] = "test_data_7111.txt";
test_data_files[7112] = "test_data_7112.txt";
test_data_files[7113] = "test_data_7113.txt";
test_data_files[7114] = "test_data_7114.txt";
test_data_files[7115] = "test_data_7115.txt";
test_data_files[7116] = "test_data_7116.txt";
test_data_files[7117] = "test_data_7117.txt";
test_data_files[7118] = "test_data_7118.txt";
test_data_files[7119] = "test_data_7119.txt";
test_data_files[7120] = "test_data_7120.txt";
test_data_files[7121] = "test_data_7121.txt";
test_data_files[7122] = "test_data_7122.txt";
test_data_files[7123] = "test_data_7123.txt";
test_data_files[7124] = "test_data_7124.txt";
test_data_files[7125] = "test_data_7125.txt";
test_data_files[7126] = "test_data_7126.txt";
test_data_files[7127] = "test_data_7127.txt";
test_data_files[7128] = "test_data_7128.txt";
test_data_files[7129] = "test_data_7129.txt";
test_data_files[7130] = "test_data_7130.txt";
test_data_files[7131] = "test_data_7131.txt";
test_data_files[7132] = "test_data_7132.txt";
test_data_files[7133] = "test_data_7133.txt";
test_data_files[7134] = "test_data_7134.txt";
test_data_files[7135] = "test_data_7135.txt";
test_data_files[7136] = "test_data_7136.txt";
test_data_files[7137] = "test_data_7137.txt";
test_data_files[7138] = "test_data_7138.txt";
test_data_files[7139] = "test_data_7139.txt";
test_data_files[7140] = "test_data_7140.txt";
test_data_files[7141] = "test_data_7141.txt";
test_data_files[7142] = "test_data_7142.txt";
test_data_files[7143] = "test_data_7143.txt";
test_data_files[7144] = "test_data_7144.txt";
test_data_files[7145] = "test_data_7145.txt";
test_data_files[7146] = "test_data_7146.txt";
test_data_files[7147] = "test_data_7147.txt";
test_data_files[7148] = "test_data_7148.txt";
test_data_files[7149] = "test_data_7149.txt";
test_data_files[7150] = "test_data_7150.txt";
test_data_files[7151] = "test_data_7151.txt";
test_data_files[7152] = "test_data_7152.txt";
test_data_files[7153] = "test_data_7153.txt";
test_data_files[7154] = "test_data_7154.txt";
test_data_files[7155] = "test_data_7155.txt";
test_data_files[7156] = "test_data_7156.txt";
test_data_files[7157] = "test_data_7157.txt";
test_data_files[7158] = "test_data_7158.txt";
test_data_files[7159] = "test_data_7159.txt";
test_data_files[7160] = "test_data_7160.txt";
test_data_files[7161] = "test_data_7161.txt";
test_data_files[7162] = "test_data_7162.txt";
test_data_files[7163] = "test_data_7163.txt";
test_data_files[7164] = "test_data_7164.txt";
test_data_files[7165] = "test_data_7165.txt";
test_data_files[7166] = "test_data_7166.txt";
test_data_files[7167] = "test_data_7167.txt";
test_data_files[7168] = "test_data_7168.txt";
test_data_files[7169] = "test_data_7169.txt";
test_data_files[7170] = "test_data_7170.txt";
test_data_files[7171] = "test_data_7171.txt";
test_data_files[7172] = "test_data_7172.txt";
test_data_files[7173] = "test_data_7173.txt";
test_data_files[7174] = "test_data_7174.txt";
test_data_files[7175] = "test_data_7175.txt";
test_data_files[7176] = "test_data_7176.txt";
test_data_files[7177] = "test_data_7177.txt";
test_data_files[7178] = "test_data_7178.txt";
test_data_files[7179] = "test_data_7179.txt";
test_data_files[7180] = "test_data_7180.txt";
test_data_files[7181] = "test_data_7181.txt";
test_data_files[7182] = "test_data_7182.txt";
test_data_files[7183] = "test_data_7183.txt";
test_data_files[7184] = "test_data_7184.txt";
test_data_files[7185] = "test_data_7185.txt";
test_data_files[7186] = "test_data_7186.txt";
test_data_files[7187] = "test_data_7187.txt";
test_data_files[7188] = "test_data_7188.txt";
test_data_files[7189] = "test_data_7189.txt";
test_data_files[7190] = "test_data_7190.txt";
test_data_files[7191] = "test_data_7191.txt";
test_data_files[7192] = "test_data_7192.txt";
test_data_files[7193] = "test_data_7193.txt";
test_data_files[7194] = "test_data_7194.txt";
test_data_files[7195] = "test_data_7195.txt";
test_data_files[7196] = "test_data_7196.txt";
test_data_files[7197] = "test_data_7197.txt";
test_data_files[7198] = "test_data_7198.txt";
test_data_files[7199] = "test_data_7199.txt";
test_data_files[7200] = "test_data_7200.txt";
test_data_files[7201] = "test_data_7201.txt";
test_data_files[7202] = "test_data_7202.txt";
test_data_files[7203] = "test_data_7203.txt";
test_data_files[7204] = "test_data_7204.txt";
test_data_files[7205] = "test_data_7205.txt";
test_data_files[7206] = "test_data_7206.txt";
test_data_files[7207] = "test_data_7207.txt";
test_data_files[7208] = "test_data_7208.txt";
test_data_files[7209] = "test_data_7209.txt";
test_data_files[7210] = "test_data_7210.txt";
test_data_files[7211] = "test_data_7211.txt";
test_data_files[7212] = "test_data_7212.txt";
test_data_files[7213] = "test_data_7213.txt";
test_data_files[7214] = "test_data_7214.txt";
test_data_files[7215] = "test_data_7215.txt";
test_data_files[7216] = "test_data_7216.txt";
test_data_files[7217] = "test_data_7217.txt";
test_data_files[7218] = "test_data_7218.txt";
test_data_files[7219] = "test_data_7219.txt";
test_data_files[7220] = "test_data_7220.txt";
test_data_files[7221] = "test_data_7221.txt";
test_data_files[7222] = "test_data_7222.txt";
test_data_files[7223] = "test_data_7223.txt";
test_data_files[7224] = "test_data_7224.txt";
test_data_files[7225] = "test_data_7225.txt";
test_data_files[7226] = "test_data_7226.txt";
test_data_files[7227] = "test_data_7227.txt";
test_data_files[7228] = "test_data_7228.txt";
test_data_files[7229] = "test_data_7229.txt";
test_data_files[7230] = "test_data_7230.txt";
test_data_files[7231] = "test_data_7231.txt";
test_data_files[7232] = "test_data_7232.txt";
test_data_files[7233] = "test_data_7233.txt";
test_data_files[7234] = "test_data_7234.txt";
test_data_files[7235] = "test_data_7235.txt";
test_data_files[7236] = "test_data_7236.txt";
test_data_files[7237] = "test_data_7237.txt";
test_data_files[7238] = "test_data_7238.txt";
test_data_files[7239] = "test_data_7239.txt";
test_data_files[7240] = "test_data_7240.txt";
test_data_files[7241] = "test_data_7241.txt";
test_data_files[7242] = "test_data_7242.txt";
test_data_files[7243] = "test_data_7243.txt";
test_data_files[7244] = "test_data_7244.txt";
test_data_files[7245] = "test_data_7245.txt";
test_data_files[7246] = "test_data_7246.txt";
test_data_files[7247] = "test_data_7247.txt";
test_data_files[7248] = "test_data_7248.txt";
test_data_files[7249] = "test_data_7249.txt";
test_data_files[7250] = "test_data_7250.txt";
test_data_files[7251] = "test_data_7251.txt";
test_data_files[7252] = "test_data_7252.txt";
test_data_files[7253] = "test_data_7253.txt";
test_data_files[7254] = "test_data_7254.txt";
test_data_files[7255] = "test_data_7255.txt";
test_data_files[7256] = "test_data_7256.txt";
test_data_files[7257] = "test_data_7257.txt";
test_data_files[7258] = "test_data_7258.txt";
test_data_files[7259] = "test_data_7259.txt";
test_data_files[7260] = "test_data_7260.txt";
test_data_files[7261] = "test_data_7261.txt";
test_data_files[7262] = "test_data_7262.txt";
test_data_files[7263] = "test_data_7263.txt";
test_data_files[7264] = "test_data_7264.txt";
test_data_files[7265] = "test_data_7265.txt";
test_data_files[7266] = "test_data_7266.txt";
test_data_files[7267] = "test_data_7267.txt";
test_data_files[7268] = "test_data_7268.txt";
test_data_files[7269] = "test_data_7269.txt";
test_data_files[7270] = "test_data_7270.txt";
test_data_files[7271] = "test_data_7271.txt";
test_data_files[7272] = "test_data_7272.txt";
test_data_files[7273] = "test_data_7273.txt";
test_data_files[7274] = "test_data_7274.txt";
test_data_files[7275] = "test_data_7275.txt";
test_data_files[7276] = "test_data_7276.txt";
test_data_files[7277] = "test_data_7277.txt";
test_data_files[7278] = "test_data_7278.txt";
test_data_files[7279] = "test_data_7279.txt";
test_data_files[7280] = "test_data_7280.txt";
test_data_files[7281] = "test_data_7281.txt";
test_data_files[7282] = "test_data_7282.txt";
test_data_files[7283] = "test_data_7283.txt";
test_data_files[7284] = "test_data_7284.txt";
test_data_files[7285] = "test_data_7285.txt";
test_data_files[7286] = "test_data_7286.txt";
test_data_files[7287] = "test_data_7287.txt";
test_data_files[7288] = "test_data_7288.txt";
test_data_files[7289] = "test_data_7289.txt";
test_data_files[7290] = "test_data_7290.txt";
test_data_files[7291] = "test_data_7291.txt";
test_data_files[7292] = "test_data_7292.txt";
test_data_files[7293] = "test_data_7293.txt";
test_data_files[7294] = "test_data_7294.txt";
test_data_files[7295] = "test_data_7295.txt";
test_data_files[7296] = "test_data_7296.txt";
test_data_files[7297] = "test_data_7297.txt";
test_data_files[7298] = "test_data_7298.txt";
test_data_files[7299] = "test_data_7299.txt";
test_data_files[7300] = "test_data_7300.txt";
test_data_files[7301] = "test_data_7301.txt";
test_data_files[7302] = "test_data_7302.txt";
test_data_files[7303] = "test_data_7303.txt";
test_data_files[7304] = "test_data_7304.txt";
test_data_files[7305] = "test_data_7305.txt";
test_data_files[7306] = "test_data_7306.txt";
test_data_files[7307] = "test_data_7307.txt";
test_data_files[7308] = "test_data_7308.txt";
test_data_files[7309] = "test_data_7309.txt";
test_data_files[7310] = "test_data_7310.txt";
test_data_files[7311] = "test_data_7311.txt";
test_data_files[7312] = "test_data_7312.txt";
test_data_files[7313] = "test_data_7313.txt";
test_data_files[7314] = "test_data_7314.txt";
test_data_files[7315] = "test_data_7315.txt";
test_data_files[7316] = "test_data_7316.txt";
test_data_files[7317] = "test_data_7317.txt";
test_data_files[7318] = "test_data_7318.txt";
test_data_files[7319] = "test_data_7319.txt";
test_data_files[7320] = "test_data_7320.txt";
test_data_files[7321] = "test_data_7321.txt";
test_data_files[7322] = "test_data_7322.txt";
test_data_files[7323] = "test_data_7323.txt";
test_data_files[7324] = "test_data_7324.txt";
test_data_files[7325] = "test_data_7325.txt";
test_data_files[7326] = "test_data_7326.txt";
test_data_files[7327] = "test_data_7327.txt";
test_data_files[7328] = "test_data_7328.txt";
test_data_files[7329] = "test_data_7329.txt";
test_data_files[7330] = "test_data_7330.txt";
test_data_files[7331] = "test_data_7331.txt";
test_data_files[7332] = "test_data_7332.txt";
test_data_files[7333] = "test_data_7333.txt";
test_data_files[7334] = "test_data_7334.txt";
test_data_files[7335] = "test_data_7335.txt";
test_data_files[7336] = "test_data_7336.txt";
test_data_files[7337] = "test_data_7337.txt";
test_data_files[7338] = "test_data_7338.txt";
test_data_files[7339] = "test_data_7339.txt";
test_data_files[7340] = "test_data_7340.txt";
test_data_files[7341] = "test_data_7341.txt";
test_data_files[7342] = "test_data_7342.txt";
test_data_files[7343] = "test_data_7343.txt";
test_data_files[7344] = "test_data_7344.txt";
test_data_files[7345] = "test_data_7345.txt";
test_data_files[7346] = "test_data_7346.txt";
test_data_files[7347] = "test_data_7347.txt";
test_data_files[7348] = "test_data_7348.txt";
test_data_files[7349] = "test_data_7349.txt";
test_data_files[7350] = "test_data_7350.txt";
test_data_files[7351] = "test_data_7351.txt";
test_data_files[7352] = "test_data_7352.txt";
test_data_files[7353] = "test_data_7353.txt";
test_data_files[7354] = "test_data_7354.txt";
test_data_files[7355] = "test_data_7355.txt";
test_data_files[7356] = "test_data_7356.txt";
test_data_files[7357] = "test_data_7357.txt";
test_data_files[7358] = "test_data_7358.txt";
test_data_files[7359] = "test_data_7359.txt";
test_data_files[7360] = "test_data_7360.txt";
test_data_files[7361] = "test_data_7361.txt";
test_data_files[7362] = "test_data_7362.txt";
test_data_files[7363] = "test_data_7363.txt";
test_data_files[7364] = "test_data_7364.txt";
test_data_files[7365] = "test_data_7365.txt";
test_data_files[7366] = "test_data_7366.txt";
test_data_files[7367] = "test_data_7367.txt";
test_data_files[7368] = "test_data_7368.txt";
test_data_files[7369] = "test_data_7369.txt";
test_data_files[7370] = "test_data_7370.txt";
test_data_files[7371] = "test_data_7371.txt";
test_data_files[7372] = "test_data_7372.txt";
test_data_files[7373] = "test_data_7373.txt";
test_data_files[7374] = "test_data_7374.txt";
test_data_files[7375] = "test_data_7375.txt";
test_data_files[7376] = "test_data_7376.txt";
test_data_files[7377] = "test_data_7377.txt";
test_data_files[7378] = "test_data_7378.txt";
test_data_files[7379] = "test_data_7379.txt";
test_data_files[7380] = "test_data_7380.txt";
test_data_files[7381] = "test_data_7381.txt";
test_data_files[7382] = "test_data_7382.txt";
test_data_files[7383] = "test_data_7383.txt";
test_data_files[7384] = "test_data_7384.txt";
test_data_files[7385] = "test_data_7385.txt";
test_data_files[7386] = "test_data_7386.txt";
test_data_files[7387] = "test_data_7387.txt";
test_data_files[7388] = "test_data_7388.txt";
test_data_files[7389] = "test_data_7389.txt";
test_data_files[7390] = "test_data_7390.txt";
test_data_files[7391] = "test_data_7391.txt";
test_data_files[7392] = "test_data_7392.txt";
test_data_files[7393] = "test_data_7393.txt";
test_data_files[7394] = "test_data_7394.txt";
test_data_files[7395] = "test_data_7395.txt";
test_data_files[7396] = "test_data_7396.txt";
test_data_files[7397] = "test_data_7397.txt";
test_data_files[7398] = "test_data_7398.txt";
test_data_files[7399] = "test_data_7399.txt";
test_data_files[7400] = "test_data_7400.txt";
test_data_files[7401] = "test_data_7401.txt";
test_data_files[7402] = "test_data_7402.txt";
test_data_files[7403] = "test_data_7403.txt";
test_data_files[7404] = "test_data_7404.txt";
test_data_files[7405] = "test_data_7405.txt";
test_data_files[7406] = "test_data_7406.txt";
test_data_files[7407] = "test_data_7407.txt";
test_data_files[7408] = "test_data_7408.txt";
test_data_files[7409] = "test_data_7409.txt";
test_data_files[7410] = "test_data_7410.txt";
test_data_files[7411] = "test_data_7411.txt";
test_data_files[7412] = "test_data_7412.txt";
test_data_files[7413] = "test_data_7413.txt";
test_data_files[7414] = "test_data_7414.txt";
test_data_files[7415] = "test_data_7415.txt";
test_data_files[7416] = "test_data_7416.txt";
test_data_files[7417] = "test_data_7417.txt";
test_data_files[7418] = "test_data_7418.txt";
test_data_files[7419] = "test_data_7419.txt";
test_data_files[7420] = "test_data_7420.txt";
test_data_files[7421] = "test_data_7421.txt";
test_data_files[7422] = "test_data_7422.txt";
test_data_files[7423] = "test_data_7423.txt";
test_data_files[7424] = "test_data_7424.txt";
test_data_files[7425] = "test_data_7425.txt";
test_data_files[7426] = "test_data_7426.txt";
test_data_files[7427] = "test_data_7427.txt";
test_data_files[7428] = "test_data_7428.txt";
test_data_files[7429] = "test_data_7429.txt";
test_data_files[7430] = "test_data_7430.txt";
test_data_files[7431] = "test_data_7431.txt";
test_data_files[7432] = "test_data_7432.txt";
test_data_files[7433] = "test_data_7433.txt";
test_data_files[7434] = "test_data_7434.txt";
test_data_files[7435] = "test_data_7435.txt";
test_data_files[7436] = "test_data_7436.txt";
test_data_files[7437] = "test_data_7437.txt";
test_data_files[7438] = "test_data_7438.txt";
test_data_files[7439] = "test_data_7439.txt";
test_data_files[7440] = "test_data_7440.txt";
test_data_files[7441] = "test_data_7441.txt";
test_data_files[7442] = "test_data_7442.txt";
test_data_files[7443] = "test_data_7443.txt";
test_data_files[7444] = "test_data_7444.txt";
test_data_files[7445] = "test_data_7445.txt";
test_data_files[7446] = "test_data_7446.txt";
test_data_files[7447] = "test_data_7447.txt";
test_data_files[7448] = "test_data_7448.txt";
test_data_files[7449] = "test_data_7449.txt";
test_data_files[7450] = "test_data_7450.txt";
test_data_files[7451] = "test_data_7451.txt";
test_data_files[7452] = "test_data_7452.txt";
test_data_files[7453] = "test_data_7453.txt";
test_data_files[7454] = "test_data_7454.txt";
test_data_files[7455] = "test_data_7455.txt";
test_data_files[7456] = "test_data_7456.txt";
test_data_files[7457] = "test_data_7457.txt";
test_data_files[7458] = "test_data_7458.txt";
test_data_files[7459] = "test_data_7459.txt";
test_data_files[7460] = "test_data_7460.txt";
test_data_files[7461] = "test_data_7461.txt";
test_data_files[7462] = "test_data_7462.txt";
test_data_files[7463] = "test_data_7463.txt";
test_data_files[7464] = "test_data_7464.txt";
test_data_files[7465] = "test_data_7465.txt";
test_data_files[7466] = "test_data_7466.txt";
test_data_files[7467] = "test_data_7467.txt";
test_data_files[7468] = "test_data_7468.txt";
test_data_files[7469] = "test_data_7469.txt";
test_data_files[7470] = "test_data_7470.txt";
test_data_files[7471] = "test_data_7471.txt";
test_data_files[7472] = "test_data_7472.txt";
test_data_files[7473] = "test_data_7473.txt";
test_data_files[7474] = "test_data_7474.txt";
test_data_files[7475] = "test_data_7475.txt";
test_data_files[7476] = "test_data_7476.txt";
test_data_files[7477] = "test_data_7477.txt";
test_data_files[7478] = "test_data_7478.txt";
test_data_files[7479] = "test_data_7479.txt";
test_data_files[7480] = "test_data_7480.txt";
test_data_files[7481] = "test_data_7481.txt";
test_data_files[7482] = "test_data_7482.txt";
test_data_files[7483] = "test_data_7483.txt";
test_data_files[7484] = "test_data_7484.txt";
test_data_files[7485] = "test_data_7485.txt";
test_data_files[7486] = "test_data_7486.txt";
test_data_files[7487] = "test_data_7487.txt";
test_data_files[7488] = "test_data_7488.txt";
test_data_files[7489] = "test_data_7489.txt";
test_data_files[7490] = "test_data_7490.txt";
test_data_files[7491] = "test_data_7491.txt";
test_data_files[7492] = "test_data_7492.txt";
test_data_files[7493] = "test_data_7493.txt";
test_data_files[7494] = "test_data_7494.txt";
test_data_files[7495] = "test_data_7495.txt";
test_data_files[7496] = "test_data_7496.txt";
test_data_files[7497] = "test_data_7497.txt";
test_data_files[7498] = "test_data_7498.txt";
test_data_files[7499] = "test_data_7499.txt";
test_data_files[7500] = "test_data_7500.txt";
test_data_files[7501] = "test_data_7501.txt";
test_data_files[7502] = "test_data_7502.txt";
test_data_files[7503] = "test_data_7503.txt";
test_data_files[7504] = "test_data_7504.txt";
test_data_files[7505] = "test_data_7505.txt";
test_data_files[7506] = "test_data_7506.txt";
test_data_files[7507] = "test_data_7507.txt";
test_data_files[7508] = "test_data_7508.txt";
test_data_files[7509] = "test_data_7509.txt";
test_data_files[7510] = "test_data_7510.txt";
test_data_files[7511] = "test_data_7511.txt";
test_data_files[7512] = "test_data_7512.txt";
test_data_files[7513] = "test_data_7513.txt";
test_data_files[7514] = "test_data_7514.txt";
test_data_files[7515] = "test_data_7515.txt";
test_data_files[7516] = "test_data_7516.txt";
test_data_files[7517] = "test_data_7517.txt";
test_data_files[7518] = "test_data_7518.txt";
test_data_files[7519] = "test_data_7519.txt";
test_data_files[7520] = "test_data_7520.txt";
test_data_files[7521] = "test_data_7521.txt";
test_data_files[7522] = "test_data_7522.txt";
test_data_files[7523] = "test_data_7523.txt";
test_data_files[7524] = "test_data_7524.txt";
test_data_files[7525] = "test_data_7525.txt";
test_data_files[7526] = "test_data_7526.txt";
test_data_files[7527] = "test_data_7527.txt";
test_data_files[7528] = "test_data_7528.txt";
test_data_files[7529] = "test_data_7529.txt";
test_data_files[7530] = "test_data_7530.txt";
test_data_files[7531] = "test_data_7531.txt";
test_data_files[7532] = "test_data_7532.txt";
test_data_files[7533] = "test_data_7533.txt";
test_data_files[7534] = "test_data_7534.txt";
test_data_files[7535] = "test_data_7535.txt";
test_data_files[7536] = "test_data_7536.txt";
test_data_files[7537] = "test_data_7537.txt";
test_data_files[7538] = "test_data_7538.txt";
test_data_files[7539] = "test_data_7539.txt";
test_data_files[7540] = "test_data_7540.txt";
test_data_files[7541] = "test_data_7541.txt";
test_data_files[7542] = "test_data_7542.txt";
test_data_files[7543] = "test_data_7543.txt";
test_data_files[7544] = "test_data_7544.txt";
test_data_files[7545] = "test_data_7545.txt";
test_data_files[7546] = "test_data_7546.txt";
test_data_files[7547] = "test_data_7547.txt";
test_data_files[7548] = "test_data_7548.txt";
test_data_files[7549] = "test_data_7549.txt";
test_data_files[7550] = "test_data_7550.txt";
test_data_files[7551] = "test_data_7551.txt";
test_data_files[7552] = "test_data_7552.txt";
test_data_files[7553] = "test_data_7553.txt";
test_data_files[7554] = "test_data_7554.txt";
test_data_files[7555] = "test_data_7555.txt";
test_data_files[7556] = "test_data_7556.txt";
test_data_files[7557] = "test_data_7557.txt";
test_data_files[7558] = "test_data_7558.txt";
test_data_files[7559] = "test_data_7559.txt";
test_data_files[7560] = "test_data_7560.txt";
test_data_files[7561] = "test_data_7561.txt";
test_data_files[7562] = "test_data_7562.txt";
test_data_files[7563] = "test_data_7563.txt";
test_data_files[7564] = "test_data_7564.txt";
test_data_files[7565] = "test_data_7565.txt";
test_data_files[7566] = "test_data_7566.txt";
test_data_files[7567] = "test_data_7567.txt";
test_data_files[7568] = "test_data_7568.txt";
test_data_files[7569] = "test_data_7569.txt";
test_data_files[7570] = "test_data_7570.txt";
test_data_files[7571] = "test_data_7571.txt";
test_data_files[7572] = "test_data_7572.txt";
test_data_files[7573] = "test_data_7573.txt";
test_data_files[7574] = "test_data_7574.txt";
test_data_files[7575] = "test_data_7575.txt";
test_data_files[7576] = "test_data_7576.txt";
test_data_files[7577] = "test_data_7577.txt";
test_data_files[7578] = "test_data_7578.txt";
test_data_files[7579] = "test_data_7579.txt";
test_data_files[7580] = "test_data_7580.txt";
test_data_files[7581] = "test_data_7581.txt";
test_data_files[7582] = "test_data_7582.txt";
test_data_files[7583] = "test_data_7583.txt";
test_data_files[7584] = "test_data_7584.txt";
test_data_files[7585] = "test_data_7585.txt";
test_data_files[7586] = "test_data_7586.txt";
test_data_files[7587] = "test_data_7587.txt";
test_data_files[7588] = "test_data_7588.txt";
test_data_files[7589] = "test_data_7589.txt";
test_data_files[7590] = "test_data_7590.txt";
test_data_files[7591] = "test_data_7591.txt";
test_data_files[7592] = "test_data_7592.txt";
test_data_files[7593] = "test_data_7593.txt";
test_data_files[7594] = "test_data_7594.txt";
test_data_files[7595] = "test_data_7595.txt";
test_data_files[7596] = "test_data_7596.txt";
test_data_files[7597] = "test_data_7597.txt";
test_data_files[7598] = "test_data_7598.txt";
test_data_files[7599] = "test_data_7599.txt";
test_data_files[7600] = "test_data_7600.txt";
test_data_files[7601] = "test_data_7601.txt";
test_data_files[7602] = "test_data_7602.txt";
test_data_files[7603] = "test_data_7603.txt";
test_data_files[7604] = "test_data_7604.txt";
test_data_files[7605] = "test_data_7605.txt";
test_data_files[7606] = "test_data_7606.txt";
test_data_files[7607] = "test_data_7607.txt";
test_data_files[7608] = "test_data_7608.txt";
test_data_files[7609] = "test_data_7609.txt";
test_data_files[7610] = "test_data_7610.txt";
test_data_files[7611] = "test_data_7611.txt";
test_data_files[7612] = "test_data_7612.txt";
test_data_files[7613] = "test_data_7613.txt";
test_data_files[7614] = "test_data_7614.txt";
test_data_files[7615] = "test_data_7615.txt";
test_data_files[7616] = "test_data_7616.txt";
test_data_files[7617] = "test_data_7617.txt";
test_data_files[7618] = "test_data_7618.txt";
test_data_files[7619] = "test_data_7619.txt";
test_data_files[7620] = "test_data_7620.txt";
test_data_files[7621] = "test_data_7621.txt";
test_data_files[7622] = "test_data_7622.txt";
test_data_files[7623] = "test_data_7623.txt";
test_data_files[7624] = "test_data_7624.txt";
test_data_files[7625] = "test_data_7625.txt";
test_data_files[7626] = "test_data_7626.txt";
test_data_files[7627] = "test_data_7627.txt";
test_data_files[7628] = "test_data_7628.txt";
test_data_files[7629] = "test_data_7629.txt";
test_data_files[7630] = "test_data_7630.txt";
test_data_files[7631] = "test_data_7631.txt";
test_data_files[7632] = "test_data_7632.txt";
test_data_files[7633] = "test_data_7633.txt";
test_data_files[7634] = "test_data_7634.txt";
test_data_files[7635] = "test_data_7635.txt";
test_data_files[7636] = "test_data_7636.txt";
test_data_files[7637] = "test_data_7637.txt";
test_data_files[7638] = "test_data_7638.txt";
test_data_files[7639] = "test_data_7639.txt";
test_data_files[7640] = "test_data_7640.txt";
test_data_files[7641] = "test_data_7641.txt";
test_data_files[7642] = "test_data_7642.txt";
test_data_files[7643] = "test_data_7643.txt";
test_data_files[7644] = "test_data_7644.txt";
test_data_files[7645] = "test_data_7645.txt";
test_data_files[7646] = "test_data_7646.txt";
test_data_files[7647] = "test_data_7647.txt";
test_data_files[7648] = "test_data_7648.txt";
test_data_files[7649] = "test_data_7649.txt";
test_data_files[7650] = "test_data_7650.txt";
test_data_files[7651] = "test_data_7651.txt";
test_data_files[7652] = "test_data_7652.txt";
test_data_files[7653] = "test_data_7653.txt";
test_data_files[7654] = "test_data_7654.txt";
test_data_files[7655] = "test_data_7655.txt";
test_data_files[7656] = "test_data_7656.txt";
test_data_files[7657] = "test_data_7657.txt";
test_data_files[7658] = "test_data_7658.txt";
test_data_files[7659] = "test_data_7659.txt";
test_data_files[7660] = "test_data_7660.txt";
test_data_files[7661] = "test_data_7661.txt";
test_data_files[7662] = "test_data_7662.txt";
test_data_files[7663] = "test_data_7663.txt";
test_data_files[7664] = "test_data_7664.txt";
test_data_files[7665] = "test_data_7665.txt";
test_data_files[7666] = "test_data_7666.txt";
test_data_files[7667] = "test_data_7667.txt";
test_data_files[7668] = "test_data_7668.txt";
test_data_files[7669] = "test_data_7669.txt";
test_data_files[7670] = "test_data_7670.txt";
test_data_files[7671] = "test_data_7671.txt";
test_data_files[7672] = "test_data_7672.txt";
test_data_files[7673] = "test_data_7673.txt";
test_data_files[7674] = "test_data_7674.txt";
test_data_files[7675] = "test_data_7675.txt";
test_data_files[7676] = "test_data_7676.txt";
test_data_files[7677] = "test_data_7677.txt";
test_data_files[7678] = "test_data_7678.txt";
test_data_files[7679] = "test_data_7679.txt";
test_data_files[7680] = "test_data_7680.txt";
test_data_files[7681] = "test_data_7681.txt";
test_data_files[7682] = "test_data_7682.txt";
test_data_files[7683] = "test_data_7683.txt";
test_data_files[7684] = "test_data_7684.txt";
test_data_files[7685] = "test_data_7685.txt";
test_data_files[7686] = "test_data_7686.txt";
test_data_files[7687] = "test_data_7687.txt";
test_data_files[7688] = "test_data_7688.txt";
test_data_files[7689] = "test_data_7689.txt";
test_data_files[7690] = "test_data_7690.txt";
test_data_files[7691] = "test_data_7691.txt";
test_data_files[7692] = "test_data_7692.txt";
test_data_files[7693] = "test_data_7693.txt";
test_data_files[7694] = "test_data_7694.txt";
test_data_files[7695] = "test_data_7695.txt";
test_data_files[7696] = "test_data_7696.txt";
test_data_files[7697] = "test_data_7697.txt";
test_data_files[7698] = "test_data_7698.txt";
test_data_files[7699] = "test_data_7699.txt";
test_data_files[7700] = "test_data_7700.txt";
test_data_files[7701] = "test_data_7701.txt";
test_data_files[7702] = "test_data_7702.txt";
test_data_files[7703] = "test_data_7703.txt";
test_data_files[7704] = "test_data_7704.txt";
test_data_files[7705] = "test_data_7705.txt";
test_data_files[7706] = "test_data_7706.txt";
test_data_files[7707] = "test_data_7707.txt";
test_data_files[7708] = "test_data_7708.txt";
test_data_files[7709] = "test_data_7709.txt";
test_data_files[7710] = "test_data_7710.txt";
test_data_files[7711] = "test_data_7711.txt";
test_data_files[7712] = "test_data_7712.txt";
test_data_files[7713] = "test_data_7713.txt";
test_data_files[7714] = "test_data_7714.txt";
test_data_files[7715] = "test_data_7715.txt";
test_data_files[7716] = "test_data_7716.txt";
test_data_files[7717] = "test_data_7717.txt";
test_data_files[7718] = "test_data_7718.txt";
test_data_files[7719] = "test_data_7719.txt";
test_data_files[7720] = "test_data_7720.txt";
test_data_files[7721] = "test_data_7721.txt";
test_data_files[7722] = "test_data_7722.txt";
test_data_files[7723] = "test_data_7723.txt";
test_data_files[7724] = "test_data_7724.txt";
test_data_files[7725] = "test_data_7725.txt";
test_data_files[7726] = "test_data_7726.txt";
test_data_files[7727] = "test_data_7727.txt";
test_data_files[7728] = "test_data_7728.txt";
test_data_files[7729] = "test_data_7729.txt";
test_data_files[7730] = "test_data_7730.txt";
test_data_files[7731] = "test_data_7731.txt";
test_data_files[7732] = "test_data_7732.txt";
test_data_files[7733] = "test_data_7733.txt";
test_data_files[7734] = "test_data_7734.txt";
test_data_files[7735] = "test_data_7735.txt";
test_data_files[7736] = "test_data_7736.txt";
test_data_files[7737] = "test_data_7737.txt";
test_data_files[7738] = "test_data_7738.txt";
test_data_files[7739] = "test_data_7739.txt";
test_data_files[7740] = "test_data_7740.txt";
test_data_files[7741] = "test_data_7741.txt";
test_data_files[7742] = "test_data_7742.txt";
test_data_files[7743] = "test_data_7743.txt";
test_data_files[7744] = "test_data_7744.txt";
test_data_files[7745] = "test_data_7745.txt";
test_data_files[7746] = "test_data_7746.txt";
test_data_files[7747] = "test_data_7747.txt";
test_data_files[7748] = "test_data_7748.txt";
test_data_files[7749] = "test_data_7749.txt";
test_data_files[7750] = "test_data_7750.txt";
test_data_files[7751] = "test_data_7751.txt";
test_data_files[7752] = "test_data_7752.txt";
test_data_files[7753] = "test_data_7753.txt";
test_data_files[7754] = "test_data_7754.txt";
test_data_files[7755] = "test_data_7755.txt";
test_data_files[7756] = "test_data_7756.txt";
test_data_files[7757] = "test_data_7757.txt";
test_data_files[7758] = "test_data_7758.txt";
test_data_files[7759] = "test_data_7759.txt";
test_data_files[7760] = "test_data_7760.txt";
test_data_files[7761] = "test_data_7761.txt";
test_data_files[7762] = "test_data_7762.txt";
test_data_files[7763] = "test_data_7763.txt";
test_data_files[7764] = "test_data_7764.txt";
test_data_files[7765] = "test_data_7765.txt";
test_data_files[7766] = "test_data_7766.txt";
test_data_files[7767] = "test_data_7767.txt";
test_data_files[7768] = "test_data_7768.txt";
test_data_files[7769] = "test_data_7769.txt";
test_data_files[7770] = "test_data_7770.txt";
test_data_files[7771] = "test_data_7771.txt";
test_data_files[7772] = "test_data_7772.txt";
test_data_files[7773] = "test_data_7773.txt";
test_data_files[7774] = "test_data_7774.txt";
test_data_files[7775] = "test_data_7775.txt";
test_data_files[7776] = "test_data_7776.txt";
test_data_files[7777] = "test_data_7777.txt";
test_data_files[7778] = "test_data_7778.txt";
test_data_files[7779] = "test_data_7779.txt";
test_data_files[7780] = "test_data_7780.txt";
test_data_files[7781] = "test_data_7781.txt";
test_data_files[7782] = "test_data_7782.txt";
test_data_files[7783] = "test_data_7783.txt";
test_data_files[7784] = "test_data_7784.txt";
test_data_files[7785] = "test_data_7785.txt";
test_data_files[7786] = "test_data_7786.txt";
test_data_files[7787] = "test_data_7787.txt";
test_data_files[7788] = "test_data_7788.txt";
test_data_files[7789] = "test_data_7789.txt";
test_data_files[7790] = "test_data_7790.txt";
test_data_files[7791] = "test_data_7791.txt";
test_data_files[7792] = "test_data_7792.txt";
test_data_files[7793] = "test_data_7793.txt";
test_data_files[7794] = "test_data_7794.txt";
test_data_files[7795] = "test_data_7795.txt";
test_data_files[7796] = "test_data_7796.txt";
test_data_files[7797] = "test_data_7797.txt";
test_data_files[7798] = "test_data_7798.txt";
test_data_files[7799] = "test_data_7799.txt";
test_data_files[7800] = "test_data_7800.txt";
test_data_files[7801] = "test_data_7801.txt";
test_data_files[7802] = "test_data_7802.txt";
test_data_files[7803] = "test_data_7803.txt";
test_data_files[7804] = "test_data_7804.txt";
test_data_files[7805] = "test_data_7805.txt";
test_data_files[7806] = "test_data_7806.txt";
test_data_files[7807] = "test_data_7807.txt";
test_data_files[7808] = "test_data_7808.txt";
test_data_files[7809] = "test_data_7809.txt";
test_data_files[7810] = "test_data_7810.txt";
test_data_files[7811] = "test_data_7811.txt";
test_data_files[7812] = "test_data_7812.txt";
test_data_files[7813] = "test_data_7813.txt";
test_data_files[7814] = "test_data_7814.txt";
test_data_files[7815] = "test_data_7815.txt";
test_data_files[7816] = "test_data_7816.txt";
test_data_files[7817] = "test_data_7817.txt";
test_data_files[7818] = "test_data_7818.txt";
test_data_files[7819] = "test_data_7819.txt";
test_data_files[7820] = "test_data_7820.txt";
test_data_files[7821] = "test_data_7821.txt";
test_data_files[7822] = "test_data_7822.txt";
test_data_files[7823] = "test_data_7823.txt";
test_data_files[7824] = "test_data_7824.txt";
test_data_files[7825] = "test_data_7825.txt";
test_data_files[7826] = "test_data_7826.txt";
test_data_files[7827] = "test_data_7827.txt";
test_data_files[7828] = "test_data_7828.txt";
test_data_files[7829] = "test_data_7829.txt";
test_data_files[7830] = "test_data_7830.txt";
test_data_files[7831] = "test_data_7831.txt";
test_data_files[7832] = "test_data_7832.txt";
test_data_files[7833] = "test_data_7833.txt";
test_data_files[7834] = "test_data_7834.txt";
test_data_files[7835] = "test_data_7835.txt";
test_data_files[7836] = "test_data_7836.txt";
test_data_files[7837] = "test_data_7837.txt";
test_data_files[7838] = "test_data_7838.txt";
test_data_files[7839] = "test_data_7839.txt";
test_data_files[7840] = "test_data_7840.txt";
test_data_files[7841] = "test_data_7841.txt";
test_data_files[7842] = "test_data_7842.txt";
test_data_files[7843] = "test_data_7843.txt";
test_data_files[7844] = "test_data_7844.txt";
test_data_files[7845] = "test_data_7845.txt";
test_data_files[7846] = "test_data_7846.txt";
test_data_files[7847] = "test_data_7847.txt";
test_data_files[7848] = "test_data_7848.txt";
test_data_files[7849] = "test_data_7849.txt";
test_data_files[7850] = "test_data_7850.txt";
test_data_files[7851] = "test_data_7851.txt";
test_data_files[7852] = "test_data_7852.txt";
test_data_files[7853] = "test_data_7853.txt";
test_data_files[7854] = "test_data_7854.txt";
test_data_files[7855] = "test_data_7855.txt";
test_data_files[7856] = "test_data_7856.txt";
test_data_files[7857] = "test_data_7857.txt";
test_data_files[7858] = "test_data_7858.txt";
test_data_files[7859] = "test_data_7859.txt";
test_data_files[7860] = "test_data_7860.txt";
test_data_files[7861] = "test_data_7861.txt";
test_data_files[7862] = "test_data_7862.txt";
test_data_files[7863] = "test_data_7863.txt";
test_data_files[7864] = "test_data_7864.txt";
test_data_files[7865] = "test_data_7865.txt";
test_data_files[7866] = "test_data_7866.txt";
test_data_files[7867] = "test_data_7867.txt";
test_data_files[7868] = "test_data_7868.txt";
test_data_files[7869] = "test_data_7869.txt";
test_data_files[7870] = "test_data_7870.txt";
test_data_files[7871] = "test_data_7871.txt";
test_data_files[7872] = "test_data_7872.txt";
test_data_files[7873] = "test_data_7873.txt";
test_data_files[7874] = "test_data_7874.txt";
test_data_files[7875] = "test_data_7875.txt";
test_data_files[7876] = "test_data_7876.txt";
test_data_files[7877] = "test_data_7877.txt";
test_data_files[7878] = "test_data_7878.txt";
test_data_files[7879] = "test_data_7879.txt";
test_data_files[7880] = "test_data_7880.txt";
test_data_files[7881] = "test_data_7881.txt";
test_data_files[7882] = "test_data_7882.txt";
test_data_files[7883] = "test_data_7883.txt";
test_data_files[7884] = "test_data_7884.txt";
test_data_files[7885] = "test_data_7885.txt";
test_data_files[7886] = "test_data_7886.txt";
test_data_files[7887] = "test_data_7887.txt";
test_data_files[7888] = "test_data_7888.txt";
test_data_files[7889] = "test_data_7889.txt";
test_data_files[7890] = "test_data_7890.txt";
test_data_files[7891] = "test_data_7891.txt";
test_data_files[7892] = "test_data_7892.txt";
test_data_files[7893] = "test_data_7893.txt";
test_data_files[7894] = "test_data_7894.txt";
test_data_files[7895] = "test_data_7895.txt";
test_data_files[7896] = "test_data_7896.txt";
test_data_files[7897] = "test_data_7897.txt";
test_data_files[7898] = "test_data_7898.txt";
test_data_files[7899] = "test_data_7899.txt";
test_data_files[7900] = "test_data_7900.txt";
test_data_files[7901] = "test_data_7901.txt";
test_data_files[7902] = "test_data_7902.txt";
test_data_files[7903] = "test_data_7903.txt";
test_data_files[7904] = "test_data_7904.txt";
test_data_files[7905] = "test_data_7905.txt";
test_data_files[7906] = "test_data_7906.txt";
test_data_files[7907] = "test_data_7907.txt";
test_data_files[7908] = "test_data_7908.txt";
test_data_files[7909] = "test_data_7909.txt";
test_data_files[7910] = "test_data_7910.txt";
test_data_files[7911] = "test_data_7911.txt";
test_data_files[7912] = "test_data_7912.txt";
test_data_files[7913] = "test_data_7913.txt";
test_data_files[7914] = "test_data_7914.txt";
test_data_files[7915] = "test_data_7915.txt";
test_data_files[7916] = "test_data_7916.txt";
test_data_files[7917] = "test_data_7917.txt";
test_data_files[7918] = "test_data_7918.txt";
test_data_files[7919] = "test_data_7919.txt";
test_data_files[7920] = "test_data_7920.txt";
test_data_files[7921] = "test_data_7921.txt";
test_data_files[7922] = "test_data_7922.txt";
test_data_files[7923] = "test_data_7923.txt";
test_data_files[7924] = "test_data_7924.txt";
test_data_files[7925] = "test_data_7925.txt";
test_data_files[7926] = "test_data_7926.txt";
test_data_files[7927] = "test_data_7927.txt";
test_data_files[7928] = "test_data_7928.txt";
test_data_files[7929] = "test_data_7929.txt";
test_data_files[7930] = "test_data_7930.txt";
test_data_files[7931] = "test_data_7931.txt";
test_data_files[7932] = "test_data_7932.txt";
test_data_files[7933] = "test_data_7933.txt";
test_data_files[7934] = "test_data_7934.txt";
test_data_files[7935] = "test_data_7935.txt";
test_data_files[7936] = "test_data_7936.txt";
test_data_files[7937] = "test_data_7937.txt";
test_data_files[7938] = "test_data_7938.txt";
test_data_files[7939] = "test_data_7939.txt";
test_data_files[7940] = "test_data_7940.txt";
test_data_files[7941] = "test_data_7941.txt";
test_data_files[7942] = "test_data_7942.txt";
test_data_files[7943] = "test_data_7943.txt";
test_data_files[7944] = "test_data_7944.txt";
test_data_files[7945] = "test_data_7945.txt";
test_data_files[7946] = "test_data_7946.txt";
test_data_files[7947] = "test_data_7947.txt";
test_data_files[7948] = "test_data_7948.txt";
test_data_files[7949] = "test_data_7949.txt";
test_data_files[7950] = "test_data_7950.txt";
test_data_files[7951] = "test_data_7951.txt";
test_data_files[7952] = "test_data_7952.txt";
test_data_files[7953] = "test_data_7953.txt";
test_data_files[7954] = "test_data_7954.txt";
test_data_files[7955] = "test_data_7955.txt";
test_data_files[7956] = "test_data_7956.txt";
test_data_files[7957] = "test_data_7957.txt";
test_data_files[7958] = "test_data_7958.txt";
test_data_files[7959] = "test_data_7959.txt";
test_data_files[7960] = "test_data_7960.txt";
test_data_files[7961] = "test_data_7961.txt";
test_data_files[7962] = "test_data_7962.txt";
test_data_files[7963] = "test_data_7963.txt";
test_data_files[7964] = "test_data_7964.txt";
test_data_files[7965] = "test_data_7965.txt";
test_data_files[7966] = "test_data_7966.txt";
test_data_files[7967] = "test_data_7967.txt";
test_data_files[7968] = "test_data_7968.txt";
test_data_files[7969] = "test_data_7969.txt";
test_data_files[7970] = "test_data_7970.txt";
test_data_files[7971] = "test_data_7971.txt";
test_data_files[7972] = "test_data_7972.txt";
test_data_files[7973] = "test_data_7973.txt";
test_data_files[7974] = "test_data_7974.txt";
test_data_files[7975] = "test_data_7975.txt";
test_data_files[7976] = "test_data_7976.txt";
test_data_files[7977] = "test_data_7977.txt";
test_data_files[7978] = "test_data_7978.txt";
test_data_files[7979] = "test_data_7979.txt";
test_data_files[7980] = "test_data_7980.txt";
test_data_files[7981] = "test_data_7981.txt";
test_data_files[7982] = "test_data_7982.txt";
test_data_files[7983] = "test_data_7983.txt";
test_data_files[7984] = "test_data_7984.txt";
test_data_files[7985] = "test_data_7985.txt";
test_data_files[7986] = "test_data_7986.txt";
test_data_files[7987] = "test_data_7987.txt";
test_data_files[7988] = "test_data_7988.txt";
test_data_files[7989] = "test_data_7989.txt";
test_data_files[7990] = "test_data_7990.txt";
test_data_files[7991] = "test_data_7991.txt";
test_data_files[7992] = "test_data_7992.txt";
test_data_files[7993] = "test_data_7993.txt";
test_data_files[7994] = "test_data_7994.txt";
test_data_files[7995] = "test_data_7995.txt";
test_data_files[7996] = "test_data_7996.txt";
test_data_files[7997] = "test_data_7997.txt";
test_data_files[7998] = "test_data_7998.txt";
test_data_files[7999] = "test_data_7999.txt";
test_data_files[8000] = "test_data_8000.txt";
test_data_files[8001] = "test_data_8001.txt";
test_data_files[8002] = "test_data_8002.txt";
test_data_files[8003] = "test_data_8003.txt";
test_data_files[8004] = "test_data_8004.txt";
test_data_files[8005] = "test_data_8005.txt";
test_data_files[8006] = "test_data_8006.txt";
test_data_files[8007] = "test_data_8007.txt";
test_data_files[8008] = "test_data_8008.txt";
test_data_files[8009] = "test_data_8009.txt";
test_data_files[8010] = "test_data_8010.txt";
test_data_files[8011] = "test_data_8011.txt";
test_data_files[8012] = "test_data_8012.txt";
test_data_files[8013] = "test_data_8013.txt";
test_data_files[8014] = "test_data_8014.txt";
test_data_files[8015] = "test_data_8015.txt";
test_data_files[8016] = "test_data_8016.txt";
test_data_files[8017] = "test_data_8017.txt";
test_data_files[8018] = "test_data_8018.txt";
test_data_files[8019] = "test_data_8019.txt";
test_data_files[8020] = "test_data_8020.txt";
test_data_files[8021] = "test_data_8021.txt";
test_data_files[8022] = "test_data_8022.txt";
test_data_files[8023] = "test_data_8023.txt";
test_data_files[8024] = "test_data_8024.txt";
test_data_files[8025] = "test_data_8025.txt";
test_data_files[8026] = "test_data_8026.txt";
test_data_files[8027] = "test_data_8027.txt";
test_data_files[8028] = "test_data_8028.txt";
test_data_files[8029] = "test_data_8029.txt";
test_data_files[8030] = "test_data_8030.txt";
test_data_files[8031] = "test_data_8031.txt";
test_data_files[8032] = "test_data_8032.txt";
test_data_files[8033] = "test_data_8033.txt";
test_data_files[8034] = "test_data_8034.txt";
test_data_files[8035] = "test_data_8035.txt";
test_data_files[8036] = "test_data_8036.txt";
test_data_files[8037] = "test_data_8037.txt";
test_data_files[8038] = "test_data_8038.txt";
test_data_files[8039] = "test_data_8039.txt";
test_data_files[8040] = "test_data_8040.txt";
test_data_files[8041] = "test_data_8041.txt";
test_data_files[8042] = "test_data_8042.txt";
test_data_files[8043] = "test_data_8043.txt";
test_data_files[8044] = "test_data_8044.txt";
test_data_files[8045] = "test_data_8045.txt";
test_data_files[8046] = "test_data_8046.txt";
test_data_files[8047] = "test_data_8047.txt";
test_data_files[8048] = "test_data_8048.txt";
test_data_files[8049] = "test_data_8049.txt";
test_data_files[8050] = "test_data_8050.txt";
test_data_files[8051] = "test_data_8051.txt";
test_data_files[8052] = "test_data_8052.txt";
test_data_files[8053] = "test_data_8053.txt";
test_data_files[8054] = "test_data_8054.txt";
test_data_files[8055] = "test_data_8055.txt";
test_data_files[8056] = "test_data_8056.txt";
test_data_files[8057] = "test_data_8057.txt";
test_data_files[8058] = "test_data_8058.txt";
test_data_files[8059] = "test_data_8059.txt";
test_data_files[8060] = "test_data_8060.txt";
test_data_files[8061] = "test_data_8061.txt";
test_data_files[8062] = "test_data_8062.txt";
test_data_files[8063] = "test_data_8063.txt";
test_data_files[8064] = "test_data_8064.txt";
test_data_files[8065] = "test_data_8065.txt";
test_data_files[8066] = "test_data_8066.txt";
test_data_files[8067] = "test_data_8067.txt";
test_data_files[8068] = "test_data_8068.txt";
test_data_files[8069] = "test_data_8069.txt";
test_data_files[8070] = "test_data_8070.txt";
test_data_files[8071] = "test_data_8071.txt";
test_data_files[8072] = "test_data_8072.txt";
test_data_files[8073] = "test_data_8073.txt";
test_data_files[8074] = "test_data_8074.txt";
test_data_files[8075] = "test_data_8075.txt";
test_data_files[8076] = "test_data_8076.txt";
test_data_files[8077] = "test_data_8077.txt";
test_data_files[8078] = "test_data_8078.txt";
test_data_files[8079] = "test_data_8079.txt";
test_data_files[8080] = "test_data_8080.txt";
test_data_files[8081] = "test_data_8081.txt";
test_data_files[8082] = "test_data_8082.txt";
test_data_files[8083] = "test_data_8083.txt";
test_data_files[8084] = "test_data_8084.txt";
test_data_files[8085] = "test_data_8085.txt";
test_data_files[8086] = "test_data_8086.txt";
test_data_files[8087] = "test_data_8087.txt";
test_data_files[8088] = "test_data_8088.txt";
test_data_files[8089] = "test_data_8089.txt";
test_data_files[8090] = "test_data_8090.txt";
test_data_files[8091] = "test_data_8091.txt";
test_data_files[8092] = "test_data_8092.txt";
test_data_files[8093] = "test_data_8093.txt";
test_data_files[8094] = "test_data_8094.txt";
test_data_files[8095] = "test_data_8095.txt";
test_data_files[8096] = "test_data_8096.txt";
test_data_files[8097] = "test_data_8097.txt";
test_data_files[8098] = "test_data_8098.txt";
test_data_files[8099] = "test_data_8099.txt";
test_data_files[8100] = "test_data_8100.txt";
test_data_files[8101] = "test_data_8101.txt";
test_data_files[8102] = "test_data_8102.txt";
test_data_files[8103] = "test_data_8103.txt";
test_data_files[8104] = "test_data_8104.txt";
test_data_files[8105] = "test_data_8105.txt";
test_data_files[8106] = "test_data_8106.txt";
test_data_files[8107] = "test_data_8107.txt";
test_data_files[8108] = "test_data_8108.txt";
test_data_files[8109] = "test_data_8109.txt";
test_data_files[8110] = "test_data_8110.txt";
test_data_files[8111] = "test_data_8111.txt";
test_data_files[8112] = "test_data_8112.txt";
test_data_files[8113] = "test_data_8113.txt";
test_data_files[8114] = "test_data_8114.txt";
test_data_files[8115] = "test_data_8115.txt";
test_data_files[8116] = "test_data_8116.txt";
test_data_files[8117] = "test_data_8117.txt";
test_data_files[8118] = "test_data_8118.txt";
test_data_files[8119] = "test_data_8119.txt";
test_data_files[8120] = "test_data_8120.txt";
test_data_files[8121] = "test_data_8121.txt";
test_data_files[8122] = "test_data_8122.txt";
test_data_files[8123] = "test_data_8123.txt";
test_data_files[8124] = "test_data_8124.txt";
test_data_files[8125] = "test_data_8125.txt";
test_data_files[8126] = "test_data_8126.txt";
test_data_files[8127] = "test_data_8127.txt";
test_data_files[8128] = "test_data_8128.txt";
test_data_files[8129] = "test_data_8129.txt";
test_data_files[8130] = "test_data_8130.txt";
test_data_files[8131] = "test_data_8131.txt";
test_data_files[8132] = "test_data_8132.txt";
test_data_files[8133] = "test_data_8133.txt";
test_data_files[8134] = "test_data_8134.txt";
test_data_files[8135] = "test_data_8135.txt";
test_data_files[8136] = "test_data_8136.txt";
test_data_files[8137] = "test_data_8137.txt";
test_data_files[8138] = "test_data_8138.txt";
test_data_files[8139] = "test_data_8139.txt";
test_data_files[8140] = "test_data_8140.txt";
test_data_files[8141] = "test_data_8141.txt";
test_data_files[8142] = "test_data_8142.txt";
test_data_files[8143] = "test_data_8143.txt";
test_data_files[8144] = "test_data_8144.txt";
test_data_files[8145] = "test_data_8145.txt";
test_data_files[8146] = "test_data_8146.txt";
test_data_files[8147] = "test_data_8147.txt";
test_data_files[8148] = "test_data_8148.txt";
test_data_files[8149] = "test_data_8149.txt";
test_data_files[8150] = "test_data_8150.txt";
test_data_files[8151] = "test_data_8151.txt";
test_data_files[8152] = "test_data_8152.txt";
test_data_files[8153] = "test_data_8153.txt";
test_data_files[8154] = "test_data_8154.txt";
test_data_files[8155] = "test_data_8155.txt";
test_data_files[8156] = "test_data_8156.txt";
test_data_files[8157] = "test_data_8157.txt";
test_data_files[8158] = "test_data_8158.txt";
test_data_files[8159] = "test_data_8159.txt";
test_data_files[8160] = "test_data_8160.txt";
test_data_files[8161] = "test_data_8161.txt";
test_data_files[8162] = "test_data_8162.txt";
test_data_files[8163] = "test_data_8163.txt";
test_data_files[8164] = "test_data_8164.txt";
test_data_files[8165] = "test_data_8165.txt";
test_data_files[8166] = "test_data_8166.txt";
test_data_files[8167] = "test_data_8167.txt";
test_data_files[8168] = "test_data_8168.txt";
test_data_files[8169] = "test_data_8169.txt";
test_data_files[8170] = "test_data_8170.txt";
test_data_files[8171] = "test_data_8171.txt";
test_data_files[8172] = "test_data_8172.txt";
test_data_files[8173] = "test_data_8173.txt";
test_data_files[8174] = "test_data_8174.txt";
test_data_files[8175] = "test_data_8175.txt";
test_data_files[8176] = "test_data_8176.txt";
test_data_files[8177] = "test_data_8177.txt";
test_data_files[8178] = "test_data_8178.txt";
test_data_files[8179] = "test_data_8179.txt";
test_data_files[8180] = "test_data_8180.txt";
test_data_files[8181] = "test_data_8181.txt";
test_data_files[8182] = "test_data_8182.txt";
test_data_files[8183] = "test_data_8183.txt";
test_data_files[8184] = "test_data_8184.txt";
test_data_files[8185] = "test_data_8185.txt";
test_data_files[8186] = "test_data_8186.txt";
test_data_files[8187] = "test_data_8187.txt";
test_data_files[8188] = "test_data_8188.txt";
test_data_files[8189] = "test_data_8189.txt";
test_data_files[8190] = "test_data_8190.txt";
test_data_files[8191] = "test_data_8191.txt";
test_data_files[8192] = "test_data_8192.txt";
test_data_files[8193] = "test_data_8193.txt";
test_data_files[8194] = "test_data_8194.txt";
test_data_files[8195] = "test_data_8195.txt";
test_data_files[8196] = "test_data_8196.txt";
test_data_files[8197] = "test_data_8197.txt";
test_data_files[8198] = "test_data_8198.txt";
test_data_files[8199] = "test_data_8199.txt";
test_data_files[8200] = "test_data_8200.txt";
test_data_files[8201] = "test_data_8201.txt";
test_data_files[8202] = "test_data_8202.txt";
test_data_files[8203] = "test_data_8203.txt";
test_data_files[8204] = "test_data_8204.txt";
test_data_files[8205] = "test_data_8205.txt";
test_data_files[8206] = "test_data_8206.txt";
test_data_files[8207] = "test_data_8207.txt";
test_data_files[8208] = "test_data_8208.txt";
test_data_files[8209] = "test_data_8209.txt";
test_data_files[8210] = "test_data_8210.txt";
test_data_files[8211] = "test_data_8211.txt";
test_data_files[8212] = "test_data_8212.txt";
test_data_files[8213] = "test_data_8213.txt";
test_data_files[8214] = "test_data_8214.txt";
test_data_files[8215] = "test_data_8215.txt";
test_data_files[8216] = "test_data_8216.txt";
test_data_files[8217] = "test_data_8217.txt";
test_data_files[8218] = "test_data_8218.txt";
test_data_files[8219] = "test_data_8219.txt";
test_data_files[8220] = "test_data_8220.txt";
test_data_files[8221] = "test_data_8221.txt";
test_data_files[8222] = "test_data_8222.txt";
test_data_files[8223] = "test_data_8223.txt";
test_data_files[8224] = "test_data_8224.txt";
test_data_files[8225] = "test_data_8225.txt";
test_data_files[8226] = "test_data_8226.txt";
test_data_files[8227] = "test_data_8227.txt";
test_data_files[8228] = "test_data_8228.txt";
test_data_files[8229] = "test_data_8229.txt";
test_data_files[8230] = "test_data_8230.txt";
test_data_files[8231] = "test_data_8231.txt";
test_data_files[8232] = "test_data_8232.txt";
test_data_files[8233] = "test_data_8233.txt";
test_data_files[8234] = "test_data_8234.txt";
test_data_files[8235] = "test_data_8235.txt";
test_data_files[8236] = "test_data_8236.txt";
test_data_files[8237] = "test_data_8237.txt";
test_data_files[8238] = "test_data_8238.txt";
test_data_files[8239] = "test_data_8239.txt";
test_data_files[8240] = "test_data_8240.txt";
test_data_files[8241] = "test_data_8241.txt";
test_data_files[8242] = "test_data_8242.txt";
test_data_files[8243] = "test_data_8243.txt";
test_data_files[8244] = "test_data_8244.txt";
test_data_files[8245] = "test_data_8245.txt";
test_data_files[8246] = "test_data_8246.txt";
test_data_files[8247] = "test_data_8247.txt";
test_data_files[8248] = "test_data_8248.txt";
test_data_files[8249] = "test_data_8249.txt";
test_data_files[8250] = "test_data_8250.txt";
test_data_files[8251] = "test_data_8251.txt";
test_data_files[8252] = "test_data_8252.txt";
test_data_files[8253] = "test_data_8253.txt";
test_data_files[8254] = "test_data_8254.txt";
test_data_files[8255] = "test_data_8255.txt";
test_data_files[8256] = "test_data_8256.txt";
test_data_files[8257] = "test_data_8257.txt";
test_data_files[8258] = "test_data_8258.txt";
test_data_files[8259] = "test_data_8259.txt";
test_data_files[8260] = "test_data_8260.txt";
test_data_files[8261] = "test_data_8261.txt";
test_data_files[8262] = "test_data_8262.txt";
test_data_files[8263] = "test_data_8263.txt";
test_data_files[8264] = "test_data_8264.txt";
test_data_files[8265] = "test_data_8265.txt";
test_data_files[8266] = "test_data_8266.txt";
test_data_files[8267] = "test_data_8267.txt";
test_data_files[8268] = "test_data_8268.txt";
test_data_files[8269] = "test_data_8269.txt";
test_data_files[8270] = "test_data_8270.txt";
test_data_files[8271] = "test_data_8271.txt";
test_data_files[8272] = "test_data_8272.txt";
test_data_files[8273] = "test_data_8273.txt";
test_data_files[8274] = "test_data_8274.txt";
test_data_files[8275] = "test_data_8275.txt";
test_data_files[8276] = "test_data_8276.txt";
test_data_files[8277] = "test_data_8277.txt";
test_data_files[8278] = "test_data_8278.txt";
test_data_files[8279] = "test_data_8279.txt";
test_data_files[8280] = "test_data_8280.txt";
test_data_files[8281] = "test_data_8281.txt";
test_data_files[8282] = "test_data_8282.txt";
test_data_files[8283] = "test_data_8283.txt";
test_data_files[8284] = "test_data_8284.txt";
test_data_files[8285] = "test_data_8285.txt";
test_data_files[8286] = "test_data_8286.txt";
test_data_files[8287] = "test_data_8287.txt";
test_data_files[8288] = "test_data_8288.txt";
test_data_files[8289] = "test_data_8289.txt";
test_data_files[8290] = "test_data_8290.txt";
test_data_files[8291] = "test_data_8291.txt";
test_data_files[8292] = "test_data_8292.txt";
test_data_files[8293] = "test_data_8293.txt";
test_data_files[8294] = "test_data_8294.txt";
test_data_files[8295] = "test_data_8295.txt";
test_data_files[8296] = "test_data_8296.txt";
test_data_files[8297] = "test_data_8297.txt";
test_data_files[8298] = "test_data_8298.txt";
test_data_files[8299] = "test_data_8299.txt";
test_data_files[8300] = "test_data_8300.txt";
test_data_files[8301] = "test_data_8301.txt";
test_data_files[8302] = "test_data_8302.txt";
test_data_files[8303] = "test_data_8303.txt";
test_data_files[8304] = "test_data_8304.txt";
test_data_files[8305] = "test_data_8305.txt";
test_data_files[8306] = "test_data_8306.txt";
test_data_files[8307] = "test_data_8307.txt";
test_data_files[8308] = "test_data_8308.txt";
test_data_files[8309] = "test_data_8309.txt";
test_data_files[8310] = "test_data_8310.txt";
test_data_files[8311] = "test_data_8311.txt";
test_data_files[8312] = "test_data_8312.txt";
test_data_files[8313] = "test_data_8313.txt";
test_data_files[8314] = "test_data_8314.txt";
test_data_files[8315] = "test_data_8315.txt";
test_data_files[8316] = "test_data_8316.txt";
test_data_files[8317] = "test_data_8317.txt";
test_data_files[8318] = "test_data_8318.txt";
test_data_files[8319] = "test_data_8319.txt";
test_data_files[8320] = "test_data_8320.txt";
test_data_files[8321] = "test_data_8321.txt";
test_data_files[8322] = "test_data_8322.txt";
test_data_files[8323] = "test_data_8323.txt";
test_data_files[8324] = "test_data_8324.txt";
test_data_files[8325] = "test_data_8325.txt";
test_data_files[8326] = "test_data_8326.txt";
test_data_files[8327] = "test_data_8327.txt";
test_data_files[8328] = "test_data_8328.txt";
test_data_files[8329] = "test_data_8329.txt";
test_data_files[8330] = "test_data_8330.txt";
test_data_files[8331] = "test_data_8331.txt";
test_data_files[8332] = "test_data_8332.txt";
test_data_files[8333] = "test_data_8333.txt";
test_data_files[8334] = "test_data_8334.txt";
test_data_files[8335] = "test_data_8335.txt";
test_data_files[8336] = "test_data_8336.txt";
test_data_files[8337] = "test_data_8337.txt";
test_data_files[8338] = "test_data_8338.txt";
test_data_files[8339] = "test_data_8339.txt";
test_data_files[8340] = "test_data_8340.txt";
test_data_files[8341] = "test_data_8341.txt";
test_data_files[8342] = "test_data_8342.txt";
test_data_files[8343] = "test_data_8343.txt";
test_data_files[8344] = "test_data_8344.txt";
test_data_files[8345] = "test_data_8345.txt";
test_data_files[8346] = "test_data_8346.txt";
test_data_files[8347] = "test_data_8347.txt";
test_data_files[8348] = "test_data_8348.txt";
test_data_files[8349] = "test_data_8349.txt";
test_data_files[8350] = "test_data_8350.txt";
test_data_files[8351] = "test_data_8351.txt";
test_data_files[8352] = "test_data_8352.txt";
test_data_files[8353] = "test_data_8353.txt";
test_data_files[8354] = "test_data_8354.txt";
test_data_files[8355] = "test_data_8355.txt";
test_data_files[8356] = "test_data_8356.txt";
test_data_files[8357] = "test_data_8357.txt";
test_data_files[8358] = "test_data_8358.txt";
test_data_files[8359] = "test_data_8359.txt";
test_data_files[8360] = "test_data_8360.txt";
test_data_files[8361] = "test_data_8361.txt";
test_data_files[8362] = "test_data_8362.txt";
test_data_files[8363] = "test_data_8363.txt";
test_data_files[8364] = "test_data_8364.txt";
test_data_files[8365] = "test_data_8365.txt";
test_data_files[8366] = "test_data_8366.txt";
test_data_files[8367] = "test_data_8367.txt";
test_data_files[8368] = "test_data_8368.txt";
test_data_files[8369] = "test_data_8369.txt";
test_data_files[8370] = "test_data_8370.txt";
test_data_files[8371] = "test_data_8371.txt";
test_data_files[8372] = "test_data_8372.txt";
test_data_files[8373] = "test_data_8373.txt";
test_data_files[8374] = "test_data_8374.txt";
test_data_files[8375] = "test_data_8375.txt";
test_data_files[8376] = "test_data_8376.txt";
test_data_files[8377] = "test_data_8377.txt";
test_data_files[8378] = "test_data_8378.txt";
test_data_files[8379] = "test_data_8379.txt";
test_data_files[8380] = "test_data_8380.txt";
test_data_files[8381] = "test_data_8381.txt";
test_data_files[8382] = "test_data_8382.txt";
test_data_files[8383] = "test_data_8383.txt";
test_data_files[8384] = "test_data_8384.txt";
test_data_files[8385] = "test_data_8385.txt";
test_data_files[8386] = "test_data_8386.txt";
test_data_files[8387] = "test_data_8387.txt";
test_data_files[8388] = "test_data_8388.txt";
test_data_files[8389] = "test_data_8389.txt";
test_data_files[8390] = "test_data_8390.txt";
test_data_files[8391] = "test_data_8391.txt";
test_data_files[8392] = "test_data_8392.txt";
test_data_files[8393] = "test_data_8393.txt";
test_data_files[8394] = "test_data_8394.txt";
test_data_files[8395] = "test_data_8395.txt";
test_data_files[8396] = "test_data_8396.txt";
test_data_files[8397] = "test_data_8397.txt";
test_data_files[8398] = "test_data_8398.txt";
test_data_files[8399] = "test_data_8399.txt";
test_data_files[8400] = "test_data_8400.txt";
test_data_files[8401] = "test_data_8401.txt";
test_data_files[8402] = "test_data_8402.txt";
test_data_files[8403] = "test_data_8403.txt";
test_data_files[8404] = "test_data_8404.txt";
test_data_files[8405] = "test_data_8405.txt";
test_data_files[8406] = "test_data_8406.txt";
test_data_files[8407] = "test_data_8407.txt";
test_data_files[8408] = "test_data_8408.txt";
test_data_files[8409] = "test_data_8409.txt";
test_data_files[8410] = "test_data_8410.txt";
test_data_files[8411] = "test_data_8411.txt";
test_data_files[8412] = "test_data_8412.txt";
test_data_files[8413] = "test_data_8413.txt";
test_data_files[8414] = "test_data_8414.txt";
test_data_files[8415] = "test_data_8415.txt";
test_data_files[8416] = "test_data_8416.txt";
test_data_files[8417] = "test_data_8417.txt";
test_data_files[8418] = "test_data_8418.txt";
test_data_files[8419] = "test_data_8419.txt";
test_data_files[8420] = "test_data_8420.txt";
test_data_files[8421] = "test_data_8421.txt";
test_data_files[8422] = "test_data_8422.txt";
test_data_files[8423] = "test_data_8423.txt";
test_data_files[8424] = "test_data_8424.txt";
test_data_files[8425] = "test_data_8425.txt";
test_data_files[8426] = "test_data_8426.txt";
test_data_files[8427] = "test_data_8427.txt";
test_data_files[8428] = "test_data_8428.txt";
test_data_files[8429] = "test_data_8429.txt";
test_data_files[8430] = "test_data_8430.txt";
test_data_files[8431] = "test_data_8431.txt";
test_data_files[8432] = "test_data_8432.txt";
test_data_files[8433] = "test_data_8433.txt";
test_data_files[8434] = "test_data_8434.txt";
test_data_files[8435] = "test_data_8435.txt";
test_data_files[8436] = "test_data_8436.txt";
test_data_files[8437] = "test_data_8437.txt";
test_data_files[8438] = "test_data_8438.txt";
test_data_files[8439] = "test_data_8439.txt";
test_data_files[8440] = "test_data_8440.txt";
test_data_files[8441] = "test_data_8441.txt";
test_data_files[8442] = "test_data_8442.txt";
test_data_files[8443] = "test_data_8443.txt";
test_data_files[8444] = "test_data_8444.txt";
test_data_files[8445] = "test_data_8445.txt";
test_data_files[8446] = "test_data_8446.txt";
test_data_files[8447] = "test_data_8447.txt";
test_data_files[8448] = "test_data_8448.txt";
test_data_files[8449] = "test_data_8449.txt";
test_data_files[8450] = "test_data_8450.txt";
test_data_files[8451] = "test_data_8451.txt";
test_data_files[8452] = "test_data_8452.txt";
test_data_files[8453] = "test_data_8453.txt";
test_data_files[8454] = "test_data_8454.txt";
test_data_files[8455] = "test_data_8455.txt";
test_data_files[8456] = "test_data_8456.txt";
test_data_files[8457] = "test_data_8457.txt";
test_data_files[8458] = "test_data_8458.txt";
test_data_files[8459] = "test_data_8459.txt";
test_data_files[8460] = "test_data_8460.txt";
test_data_files[8461] = "test_data_8461.txt";
test_data_files[8462] = "test_data_8462.txt";
test_data_files[8463] = "test_data_8463.txt";
test_data_files[8464] = "test_data_8464.txt";
test_data_files[8465] = "test_data_8465.txt";
test_data_files[8466] = "test_data_8466.txt";
test_data_files[8467] = "test_data_8467.txt";
test_data_files[8468] = "test_data_8468.txt";
test_data_files[8469] = "test_data_8469.txt";
test_data_files[8470] = "test_data_8470.txt";
test_data_files[8471] = "test_data_8471.txt";
test_data_files[8472] = "test_data_8472.txt";
test_data_files[8473] = "test_data_8473.txt";
test_data_files[8474] = "test_data_8474.txt";
test_data_files[8475] = "test_data_8475.txt";
test_data_files[8476] = "test_data_8476.txt";
test_data_files[8477] = "test_data_8477.txt";
test_data_files[8478] = "test_data_8478.txt";
test_data_files[8479] = "test_data_8479.txt";
test_data_files[8480] = "test_data_8480.txt";
test_data_files[8481] = "test_data_8481.txt";
test_data_files[8482] = "test_data_8482.txt";
test_data_files[8483] = "test_data_8483.txt";
test_data_files[8484] = "test_data_8484.txt";
test_data_files[8485] = "test_data_8485.txt";
test_data_files[8486] = "test_data_8486.txt";
test_data_files[8487] = "test_data_8487.txt";
test_data_files[8488] = "test_data_8488.txt";
test_data_files[8489] = "test_data_8489.txt";
test_data_files[8490] = "test_data_8490.txt";
test_data_files[8491] = "test_data_8491.txt";
test_data_files[8492] = "test_data_8492.txt";
test_data_files[8493] = "test_data_8493.txt";
test_data_files[8494] = "test_data_8494.txt";
test_data_files[8495] = "test_data_8495.txt";
test_data_files[8496] = "test_data_8496.txt";
test_data_files[8497] = "test_data_8497.txt";
test_data_files[8498] = "test_data_8498.txt";
test_data_files[8499] = "test_data_8499.txt";
test_data_files[8500] = "test_data_8500.txt";
test_data_files[8501] = "test_data_8501.txt";
test_data_files[8502] = "test_data_8502.txt";
test_data_files[8503] = "test_data_8503.txt";
test_data_files[8504] = "test_data_8504.txt";
test_data_files[8505] = "test_data_8505.txt";
test_data_files[8506] = "test_data_8506.txt";
test_data_files[8507] = "test_data_8507.txt";
test_data_files[8508] = "test_data_8508.txt";
test_data_files[8509] = "test_data_8509.txt";
test_data_files[8510] = "test_data_8510.txt";
test_data_files[8511] = "test_data_8511.txt";
test_data_files[8512] = "test_data_8512.txt";
test_data_files[8513] = "test_data_8513.txt";
test_data_files[8514] = "test_data_8514.txt";
test_data_files[8515] = "test_data_8515.txt";
test_data_files[8516] = "test_data_8516.txt";
test_data_files[8517] = "test_data_8517.txt";
test_data_files[8518] = "test_data_8518.txt";
test_data_files[8519] = "test_data_8519.txt";
test_data_files[8520] = "test_data_8520.txt";
test_data_files[8521] = "test_data_8521.txt";
test_data_files[8522] = "test_data_8522.txt";
test_data_files[8523] = "test_data_8523.txt";
test_data_files[8524] = "test_data_8524.txt";
test_data_files[8525] = "test_data_8525.txt";
test_data_files[8526] = "test_data_8526.txt";
test_data_files[8527] = "test_data_8527.txt";
test_data_files[8528] = "test_data_8528.txt";
test_data_files[8529] = "test_data_8529.txt";
test_data_files[8530] = "test_data_8530.txt";
test_data_files[8531] = "test_data_8531.txt";
test_data_files[8532] = "test_data_8532.txt";
test_data_files[8533] = "test_data_8533.txt";
test_data_files[8534] = "test_data_8534.txt";
test_data_files[8535] = "test_data_8535.txt";
test_data_files[8536] = "test_data_8536.txt";
test_data_files[8537] = "test_data_8537.txt";
test_data_files[8538] = "test_data_8538.txt";
test_data_files[8539] = "test_data_8539.txt";
test_data_files[8540] = "test_data_8540.txt";
test_data_files[8541] = "test_data_8541.txt";
test_data_files[8542] = "test_data_8542.txt";
test_data_files[8543] = "test_data_8543.txt";
test_data_files[8544] = "test_data_8544.txt";
test_data_files[8545] = "test_data_8545.txt";
test_data_files[8546] = "test_data_8546.txt";
test_data_files[8547] = "test_data_8547.txt";
test_data_files[8548] = "test_data_8548.txt";
test_data_files[8549] = "test_data_8549.txt";
test_data_files[8550] = "test_data_8550.txt";
test_data_files[8551] = "test_data_8551.txt";
test_data_files[8552] = "test_data_8552.txt";
test_data_files[8553] = "test_data_8553.txt";
test_data_files[8554] = "test_data_8554.txt";
test_data_files[8555] = "test_data_8555.txt";
test_data_files[8556] = "test_data_8556.txt";
test_data_files[8557] = "test_data_8557.txt";
test_data_files[8558] = "test_data_8558.txt";
test_data_files[8559] = "test_data_8559.txt";
test_data_files[8560] = "test_data_8560.txt";
test_data_files[8561] = "test_data_8561.txt";
test_data_files[8562] = "test_data_8562.txt";
test_data_files[8563] = "test_data_8563.txt";
test_data_files[8564] = "test_data_8564.txt";
test_data_files[8565] = "test_data_8565.txt";
test_data_files[8566] = "test_data_8566.txt";
test_data_files[8567] = "test_data_8567.txt";
test_data_files[8568] = "test_data_8568.txt";
test_data_files[8569] = "test_data_8569.txt";
test_data_files[8570] = "test_data_8570.txt";
test_data_files[8571] = "test_data_8571.txt";
test_data_files[8572] = "test_data_8572.txt";
test_data_files[8573] = "test_data_8573.txt";
test_data_files[8574] = "test_data_8574.txt";
test_data_files[8575] = "test_data_8575.txt";
test_data_files[8576] = "test_data_8576.txt";
test_data_files[8577] = "test_data_8577.txt";
test_data_files[8578] = "test_data_8578.txt";
test_data_files[8579] = "test_data_8579.txt";
test_data_files[8580] = "test_data_8580.txt";
test_data_files[8581] = "test_data_8581.txt";
test_data_files[8582] = "test_data_8582.txt";
test_data_files[8583] = "test_data_8583.txt";
test_data_files[8584] = "test_data_8584.txt";
test_data_files[8585] = "test_data_8585.txt";
test_data_files[8586] = "test_data_8586.txt";
test_data_files[8587] = "test_data_8587.txt";
test_data_files[8588] = "test_data_8588.txt";
test_data_files[8589] = "test_data_8589.txt";
test_data_files[8590] = "test_data_8590.txt";
test_data_files[8591] = "test_data_8591.txt";
test_data_files[8592] = "test_data_8592.txt";
test_data_files[8593] = "test_data_8593.txt";
test_data_files[8594] = "test_data_8594.txt";
test_data_files[8595] = "test_data_8595.txt";
test_data_files[8596] = "test_data_8596.txt";
test_data_files[8597] = "test_data_8597.txt";
test_data_files[8598] = "test_data_8598.txt";
test_data_files[8599] = "test_data_8599.txt";
test_data_files[8600] = "test_data_8600.txt";
test_data_files[8601] = "test_data_8601.txt";
test_data_files[8602] = "test_data_8602.txt";
test_data_files[8603] = "test_data_8603.txt";
test_data_files[8604] = "test_data_8604.txt";
test_data_files[8605] = "test_data_8605.txt";
test_data_files[8606] = "test_data_8606.txt";
test_data_files[8607] = "test_data_8607.txt";
test_data_files[8608] = "test_data_8608.txt";
test_data_files[8609] = "test_data_8609.txt";
test_data_files[8610] = "test_data_8610.txt";
test_data_files[8611] = "test_data_8611.txt";
test_data_files[8612] = "test_data_8612.txt";
test_data_files[8613] = "test_data_8613.txt";
test_data_files[8614] = "test_data_8614.txt";
test_data_files[8615] = "test_data_8615.txt";
test_data_files[8616] = "test_data_8616.txt";
test_data_files[8617] = "test_data_8617.txt";
test_data_files[8618] = "test_data_8618.txt";
test_data_files[8619] = "test_data_8619.txt";
test_data_files[8620] = "test_data_8620.txt";
test_data_files[8621] = "test_data_8621.txt";
test_data_files[8622] = "test_data_8622.txt";
test_data_files[8623] = "test_data_8623.txt";
test_data_files[8624] = "test_data_8624.txt";
test_data_files[8625] = "test_data_8625.txt";
test_data_files[8626] = "test_data_8626.txt";
test_data_files[8627] = "test_data_8627.txt";
test_data_files[8628] = "test_data_8628.txt";
test_data_files[8629] = "test_data_8629.txt";
test_data_files[8630] = "test_data_8630.txt";
test_data_files[8631] = "test_data_8631.txt";
test_data_files[8632] = "test_data_8632.txt";
test_data_files[8633] = "test_data_8633.txt";
test_data_files[8634] = "test_data_8634.txt";
test_data_files[8635] = "test_data_8635.txt";
test_data_files[8636] = "test_data_8636.txt";
test_data_files[8637] = "test_data_8637.txt";
test_data_files[8638] = "test_data_8638.txt";
test_data_files[8639] = "test_data_8639.txt";
test_data_files[8640] = "test_data_8640.txt";
test_data_files[8641] = "test_data_8641.txt";
test_data_files[8642] = "test_data_8642.txt";
test_data_files[8643] = "test_data_8643.txt";
test_data_files[8644] = "test_data_8644.txt";
test_data_files[8645] = "test_data_8645.txt";
test_data_files[8646] = "test_data_8646.txt";
test_data_files[8647] = "test_data_8647.txt";
test_data_files[8648] = "test_data_8648.txt";
test_data_files[8649] = "test_data_8649.txt";
test_data_files[8650] = "test_data_8650.txt";
test_data_files[8651] = "test_data_8651.txt";
test_data_files[8652] = "test_data_8652.txt";
test_data_files[8653] = "test_data_8653.txt";
test_data_files[8654] = "test_data_8654.txt";
test_data_files[8655] = "test_data_8655.txt";
test_data_files[8656] = "test_data_8656.txt";
test_data_files[8657] = "test_data_8657.txt";
test_data_files[8658] = "test_data_8658.txt";
test_data_files[8659] = "test_data_8659.txt";
test_data_files[8660] = "test_data_8660.txt";
test_data_files[8661] = "test_data_8661.txt";
test_data_files[8662] = "test_data_8662.txt";
test_data_files[8663] = "test_data_8663.txt";
test_data_files[8664] = "test_data_8664.txt";
test_data_files[8665] = "test_data_8665.txt";
test_data_files[8666] = "test_data_8666.txt";
test_data_files[8667] = "test_data_8667.txt";
test_data_files[8668] = "test_data_8668.txt";
test_data_files[8669] = "test_data_8669.txt";
test_data_files[8670] = "test_data_8670.txt";
test_data_files[8671] = "test_data_8671.txt";
test_data_files[8672] = "test_data_8672.txt";
test_data_files[8673] = "test_data_8673.txt";
test_data_files[8674] = "test_data_8674.txt";
test_data_files[8675] = "test_data_8675.txt";
test_data_files[8676] = "test_data_8676.txt";
test_data_files[8677] = "test_data_8677.txt";
test_data_files[8678] = "test_data_8678.txt";
test_data_files[8679] = "test_data_8679.txt";
test_data_files[8680] = "test_data_8680.txt";
test_data_files[8681] = "test_data_8681.txt";
test_data_files[8682] = "test_data_8682.txt";
test_data_files[8683] = "test_data_8683.txt";
test_data_files[8684] = "test_data_8684.txt";
test_data_files[8685] = "test_data_8685.txt";
test_data_files[8686] = "test_data_8686.txt";
test_data_files[8687] = "test_data_8687.txt";
test_data_files[8688] = "test_data_8688.txt";
test_data_files[8689] = "test_data_8689.txt";
test_data_files[8690] = "test_data_8690.txt";
test_data_files[8691] = "test_data_8691.txt";
test_data_files[8692] = "test_data_8692.txt";
test_data_files[8693] = "test_data_8693.txt";
test_data_files[8694] = "test_data_8694.txt";
test_data_files[8695] = "test_data_8695.txt";
test_data_files[8696] = "test_data_8696.txt";
test_data_files[8697] = "test_data_8697.txt";
test_data_files[8698] = "test_data_8698.txt";
test_data_files[8699] = "test_data_8699.txt";
test_data_files[8700] = "test_data_8700.txt";
test_data_files[8701] = "test_data_8701.txt";
test_data_files[8702] = "test_data_8702.txt";
test_data_files[8703] = "test_data_8703.txt";
test_data_files[8704] = "test_data_8704.txt";
test_data_files[8705] = "test_data_8705.txt";
test_data_files[8706] = "test_data_8706.txt";
test_data_files[8707] = "test_data_8707.txt";
test_data_files[8708] = "test_data_8708.txt";
test_data_files[8709] = "test_data_8709.txt";
test_data_files[8710] = "test_data_8710.txt";
test_data_files[8711] = "test_data_8711.txt";
test_data_files[8712] = "test_data_8712.txt";
test_data_files[8713] = "test_data_8713.txt";
test_data_files[8714] = "test_data_8714.txt";
test_data_files[8715] = "test_data_8715.txt";
test_data_files[8716] = "test_data_8716.txt";
test_data_files[8717] = "test_data_8717.txt";
test_data_files[8718] = "test_data_8718.txt";
test_data_files[8719] = "test_data_8719.txt";
test_data_files[8720] = "test_data_8720.txt";
test_data_files[8721] = "test_data_8721.txt";
test_data_files[8722] = "test_data_8722.txt";
test_data_files[8723] = "test_data_8723.txt";
test_data_files[8724] = "test_data_8724.txt";
test_data_files[8725] = "test_data_8725.txt";
test_data_files[8726] = "test_data_8726.txt";
test_data_files[8727] = "test_data_8727.txt";
test_data_files[8728] = "test_data_8728.txt";
test_data_files[8729] = "test_data_8729.txt";
test_data_files[8730] = "test_data_8730.txt";
test_data_files[8731] = "test_data_8731.txt";
test_data_files[8732] = "test_data_8732.txt";
test_data_files[8733] = "test_data_8733.txt";
test_data_files[8734] = "test_data_8734.txt";
test_data_files[8735] = "test_data_8735.txt";
test_data_files[8736] = "test_data_8736.txt";
test_data_files[8737] = "test_data_8737.txt";
test_data_files[8738] = "test_data_8738.txt";
test_data_files[8739] = "test_data_8739.txt";
test_data_files[8740] = "test_data_8740.txt";
test_data_files[8741] = "test_data_8741.txt";
test_data_files[8742] = "test_data_8742.txt";
test_data_files[8743] = "test_data_8743.txt";
test_data_files[8744] = "test_data_8744.txt";
test_data_files[8745] = "test_data_8745.txt";
test_data_files[8746] = "test_data_8746.txt";
test_data_files[8747] = "test_data_8747.txt";
test_data_files[8748] = "test_data_8748.txt";
test_data_files[8749] = "test_data_8749.txt";
test_data_files[8750] = "test_data_8750.txt";
test_data_files[8751] = "test_data_8751.txt";
test_data_files[8752] = "test_data_8752.txt";
test_data_files[8753] = "test_data_8753.txt";
test_data_files[8754] = "test_data_8754.txt";
test_data_files[8755] = "test_data_8755.txt";
test_data_files[8756] = "test_data_8756.txt";
test_data_files[8757] = "test_data_8757.txt";
test_data_files[8758] = "test_data_8758.txt";
test_data_files[8759] = "test_data_8759.txt";
test_data_files[8760] = "test_data_8760.txt";
test_data_files[8761] = "test_data_8761.txt";
test_data_files[8762] = "test_data_8762.txt";
test_data_files[8763] = "test_data_8763.txt";
test_data_files[8764] = "test_data_8764.txt";
test_data_files[8765] = "test_data_8765.txt";
test_data_files[8766] = "test_data_8766.txt";
test_data_files[8767] = "test_data_8767.txt";
test_data_files[8768] = "test_data_8768.txt";
test_data_files[8769] = "test_data_8769.txt";
test_data_files[8770] = "test_data_8770.txt";
test_data_files[8771] = "test_data_8771.txt";
test_data_files[8772] = "test_data_8772.txt";
test_data_files[8773] = "test_data_8773.txt";
test_data_files[8774] = "test_data_8774.txt";
test_data_files[8775] = "test_data_8775.txt";
test_data_files[8776] = "test_data_8776.txt";
test_data_files[8777] = "test_data_8777.txt";
test_data_files[8778] = "test_data_8778.txt";
test_data_files[8779] = "test_data_8779.txt";
test_data_files[8780] = "test_data_8780.txt";
test_data_files[8781] = "test_data_8781.txt";
test_data_files[8782] = "test_data_8782.txt";
test_data_files[8783] = "test_data_8783.txt";
test_data_files[8784] = "test_data_8784.txt";
test_data_files[8785] = "test_data_8785.txt";
test_data_files[8786] = "test_data_8786.txt";
test_data_files[8787] = "test_data_8787.txt";
test_data_files[8788] = "test_data_8788.txt";
test_data_files[8789] = "test_data_8789.txt";
test_data_files[8790] = "test_data_8790.txt";
test_data_files[8791] = "test_data_8791.txt";
test_data_files[8792] = "test_data_8792.txt";
test_data_files[8793] = "test_data_8793.txt";
test_data_files[8794] = "test_data_8794.txt";
test_data_files[8795] = "test_data_8795.txt";
test_data_files[8796] = "test_data_8796.txt";
test_data_files[8797] = "test_data_8797.txt";
test_data_files[8798] = "test_data_8798.txt";
test_data_files[8799] = "test_data_8799.txt";
test_data_files[8800] = "test_data_8800.txt";
test_data_files[8801] = "test_data_8801.txt";
test_data_files[8802] = "test_data_8802.txt";
test_data_files[8803] = "test_data_8803.txt";
test_data_files[8804] = "test_data_8804.txt";
test_data_files[8805] = "test_data_8805.txt";
test_data_files[8806] = "test_data_8806.txt";
test_data_files[8807] = "test_data_8807.txt";
test_data_files[8808] = "test_data_8808.txt";
test_data_files[8809] = "test_data_8809.txt";
test_data_files[8810] = "test_data_8810.txt";
test_data_files[8811] = "test_data_8811.txt";
test_data_files[8812] = "test_data_8812.txt";
test_data_files[8813] = "test_data_8813.txt";
test_data_files[8814] = "test_data_8814.txt";
test_data_files[8815] = "test_data_8815.txt";
test_data_files[8816] = "test_data_8816.txt";
test_data_files[8817] = "test_data_8817.txt";
test_data_files[8818] = "test_data_8818.txt";
test_data_files[8819] = "test_data_8819.txt";
test_data_files[8820] = "test_data_8820.txt";
test_data_files[8821] = "test_data_8821.txt";
test_data_files[8822] = "test_data_8822.txt";
test_data_files[8823] = "test_data_8823.txt";
test_data_files[8824] = "test_data_8824.txt";
test_data_files[8825] = "test_data_8825.txt";
test_data_files[8826] = "test_data_8826.txt";
test_data_files[8827] = "test_data_8827.txt";
test_data_files[8828] = "test_data_8828.txt";
test_data_files[8829] = "test_data_8829.txt";
test_data_files[8830] = "test_data_8830.txt";
test_data_files[8831] = "test_data_8831.txt";
test_data_files[8832] = "test_data_8832.txt";
test_data_files[8833] = "test_data_8833.txt";
test_data_files[8834] = "test_data_8834.txt";
test_data_files[8835] = "test_data_8835.txt";
test_data_files[8836] = "test_data_8836.txt";
test_data_files[8837] = "test_data_8837.txt";
test_data_files[8838] = "test_data_8838.txt";
test_data_files[8839] = "test_data_8839.txt";
test_data_files[8840] = "test_data_8840.txt";
test_data_files[8841] = "test_data_8841.txt";
test_data_files[8842] = "test_data_8842.txt";
test_data_files[8843] = "test_data_8843.txt";
test_data_files[8844] = "test_data_8844.txt";
test_data_files[8845] = "test_data_8845.txt";
test_data_files[8846] = "test_data_8846.txt";
test_data_files[8847] = "test_data_8847.txt";
test_data_files[8848] = "test_data_8848.txt";
test_data_files[8849] = "test_data_8849.txt";
test_data_files[8850] = "test_data_8850.txt";
test_data_files[8851] = "test_data_8851.txt";
test_data_files[8852] = "test_data_8852.txt";
test_data_files[8853] = "test_data_8853.txt";
test_data_files[8854] = "test_data_8854.txt";
test_data_files[8855] = "test_data_8855.txt";
test_data_files[8856] = "test_data_8856.txt";
test_data_files[8857] = "test_data_8857.txt";
test_data_files[8858] = "test_data_8858.txt";
test_data_files[8859] = "test_data_8859.txt";
test_data_files[8860] = "test_data_8860.txt";
test_data_files[8861] = "test_data_8861.txt";
test_data_files[8862] = "test_data_8862.txt";
test_data_files[8863] = "test_data_8863.txt";
test_data_files[8864] = "test_data_8864.txt";
test_data_files[8865] = "test_data_8865.txt";
test_data_files[8866] = "test_data_8866.txt";
test_data_files[8867] = "test_data_8867.txt";
test_data_files[8868] = "test_data_8868.txt";
test_data_files[8869] = "test_data_8869.txt";
test_data_files[8870] = "test_data_8870.txt";
test_data_files[8871] = "test_data_8871.txt";
test_data_files[8872] = "test_data_8872.txt";
test_data_files[8873] = "test_data_8873.txt";
test_data_files[8874] = "test_data_8874.txt";
test_data_files[8875] = "test_data_8875.txt";
test_data_files[8876] = "test_data_8876.txt";
test_data_files[8877] = "test_data_8877.txt";
test_data_files[8878] = "test_data_8878.txt";
test_data_files[8879] = "test_data_8879.txt";
test_data_files[8880] = "test_data_8880.txt";
test_data_files[8881] = "test_data_8881.txt";
test_data_files[8882] = "test_data_8882.txt";
test_data_files[8883] = "test_data_8883.txt";
test_data_files[8884] = "test_data_8884.txt";
test_data_files[8885] = "test_data_8885.txt";
test_data_files[8886] = "test_data_8886.txt";
test_data_files[8887] = "test_data_8887.txt";
test_data_files[8888] = "test_data_8888.txt";
test_data_files[8889] = "test_data_8889.txt";
test_data_files[8890] = "test_data_8890.txt";
test_data_files[8891] = "test_data_8891.txt";
test_data_files[8892] = "test_data_8892.txt";
test_data_files[8893] = "test_data_8893.txt";
test_data_files[8894] = "test_data_8894.txt";
test_data_files[8895] = "test_data_8895.txt";
test_data_files[8896] = "test_data_8896.txt";
test_data_files[8897] = "test_data_8897.txt";
test_data_files[8898] = "test_data_8898.txt";
test_data_files[8899] = "test_data_8899.txt";
test_data_files[8900] = "test_data_8900.txt";
test_data_files[8901] = "test_data_8901.txt";
test_data_files[8902] = "test_data_8902.txt";
test_data_files[8903] = "test_data_8903.txt";
test_data_files[8904] = "test_data_8904.txt";
test_data_files[8905] = "test_data_8905.txt";
test_data_files[8906] = "test_data_8906.txt";
test_data_files[8907] = "test_data_8907.txt";
test_data_files[8908] = "test_data_8908.txt";
test_data_files[8909] = "test_data_8909.txt";
test_data_files[8910] = "test_data_8910.txt";
test_data_files[8911] = "test_data_8911.txt";
test_data_files[8912] = "test_data_8912.txt";
test_data_files[8913] = "test_data_8913.txt";
test_data_files[8914] = "test_data_8914.txt";
test_data_files[8915] = "test_data_8915.txt";
test_data_files[8916] = "test_data_8916.txt";
test_data_files[8917] = "test_data_8917.txt";
test_data_files[8918] = "test_data_8918.txt";
test_data_files[8919] = "test_data_8919.txt";
test_data_files[8920] = "test_data_8920.txt";
test_data_files[8921] = "test_data_8921.txt";
test_data_files[8922] = "test_data_8922.txt";
test_data_files[8923] = "test_data_8923.txt";
test_data_files[8924] = "test_data_8924.txt";
test_data_files[8925] = "test_data_8925.txt";
test_data_files[8926] = "test_data_8926.txt";
test_data_files[8927] = "test_data_8927.txt";
test_data_files[8928] = "test_data_8928.txt";
test_data_files[8929] = "test_data_8929.txt";
test_data_files[8930] = "test_data_8930.txt";
test_data_files[8931] = "test_data_8931.txt";
test_data_files[8932] = "test_data_8932.txt";
test_data_files[8933] = "test_data_8933.txt";
test_data_files[8934] = "test_data_8934.txt";
test_data_files[8935] = "test_data_8935.txt";
test_data_files[8936] = "test_data_8936.txt";
test_data_files[8937] = "test_data_8937.txt";
test_data_files[8938] = "test_data_8938.txt";
test_data_files[8939] = "test_data_8939.txt";
test_data_files[8940] = "test_data_8940.txt";
test_data_files[8941] = "test_data_8941.txt";
test_data_files[8942] = "test_data_8942.txt";
test_data_files[8943] = "test_data_8943.txt";
test_data_files[8944] = "test_data_8944.txt";
test_data_files[8945] = "test_data_8945.txt";
test_data_files[8946] = "test_data_8946.txt";
test_data_files[8947] = "test_data_8947.txt";
test_data_files[8948] = "test_data_8948.txt";
test_data_files[8949] = "test_data_8949.txt";
test_data_files[8950] = "test_data_8950.txt";
test_data_files[8951] = "test_data_8951.txt";
test_data_files[8952] = "test_data_8952.txt";
test_data_files[8953] = "test_data_8953.txt";
test_data_files[8954] = "test_data_8954.txt";
test_data_files[8955] = "test_data_8955.txt";
test_data_files[8956] = "test_data_8956.txt";
test_data_files[8957] = "test_data_8957.txt";
test_data_files[8958] = "test_data_8958.txt";
test_data_files[8959] = "test_data_8959.txt";
test_data_files[8960] = "test_data_8960.txt";
test_data_files[8961] = "test_data_8961.txt";
test_data_files[8962] = "test_data_8962.txt";
test_data_files[8963] = "test_data_8963.txt";
test_data_files[8964] = "test_data_8964.txt";
test_data_files[8965] = "test_data_8965.txt";
test_data_files[8966] = "test_data_8966.txt";
test_data_files[8967] = "test_data_8967.txt";
test_data_files[8968] = "test_data_8968.txt";
test_data_files[8969] = "test_data_8969.txt";
test_data_files[8970] = "test_data_8970.txt";
test_data_files[8971] = "test_data_8971.txt";
test_data_files[8972] = "test_data_8972.txt";
test_data_files[8973] = "test_data_8973.txt";
test_data_files[8974] = "test_data_8974.txt";
test_data_files[8975] = "test_data_8975.txt";
test_data_files[8976] = "test_data_8976.txt";
test_data_files[8977] = "test_data_8977.txt";
test_data_files[8978] = "test_data_8978.txt";
test_data_files[8979] = "test_data_8979.txt";
test_data_files[8980] = "test_data_8980.txt";
test_data_files[8981] = "test_data_8981.txt";
test_data_files[8982] = "test_data_8982.txt";
test_data_files[8983] = "test_data_8983.txt";
test_data_files[8984] = "test_data_8984.txt";
test_data_files[8985] = "test_data_8985.txt";
test_data_files[8986] = "test_data_8986.txt";
test_data_files[8987] = "test_data_8987.txt";
test_data_files[8988] = "test_data_8988.txt";
test_data_files[8989] = "test_data_8989.txt";
test_data_files[8990] = "test_data_8990.txt";
test_data_files[8991] = "test_data_8991.txt";
test_data_files[8992] = "test_data_8992.txt";
test_data_files[8993] = "test_data_8993.txt";
test_data_files[8994] = "test_data_8994.txt";
test_data_files[8995] = "test_data_8995.txt";
test_data_files[8996] = "test_data_8996.txt";
test_data_files[8997] = "test_data_8997.txt";
test_data_files[8998] = "test_data_8998.txt";
test_data_files[8999] = "test_data_8999.txt";
test_data_files[9000] = "test_data_9000.txt";
test_data_files[9001] = "test_data_9001.txt";
test_data_files[9002] = "test_data_9002.txt";
test_data_files[9003] = "test_data_9003.txt";
test_data_files[9004] = "test_data_9004.txt";
test_data_files[9005] = "test_data_9005.txt";
test_data_files[9006] = "test_data_9006.txt";
test_data_files[9007] = "test_data_9007.txt";
test_data_files[9008] = "test_data_9008.txt";
test_data_files[9009] = "test_data_9009.txt";
test_data_files[9010] = "test_data_9010.txt";
test_data_files[9011] = "test_data_9011.txt";
test_data_files[9012] = "test_data_9012.txt";
test_data_files[9013] = "test_data_9013.txt";
test_data_files[9014] = "test_data_9014.txt";
test_data_files[9015] = "test_data_9015.txt";
test_data_files[9016] = "test_data_9016.txt";
test_data_files[9017] = "test_data_9017.txt";
test_data_files[9018] = "test_data_9018.txt";
test_data_files[9019] = "test_data_9019.txt";
test_data_files[9020] = "test_data_9020.txt";
test_data_files[9021] = "test_data_9021.txt";
test_data_files[9022] = "test_data_9022.txt";
test_data_files[9023] = "test_data_9023.txt";
test_data_files[9024] = "test_data_9024.txt";
test_data_files[9025] = "test_data_9025.txt";
test_data_files[9026] = "test_data_9026.txt";
test_data_files[9027] = "test_data_9027.txt";
test_data_files[9028] = "test_data_9028.txt";
test_data_files[9029] = "test_data_9029.txt";
test_data_files[9030] = "test_data_9030.txt";
test_data_files[9031] = "test_data_9031.txt";
test_data_files[9032] = "test_data_9032.txt";
test_data_files[9033] = "test_data_9033.txt";
test_data_files[9034] = "test_data_9034.txt";
test_data_files[9035] = "test_data_9035.txt";
test_data_files[9036] = "test_data_9036.txt";
test_data_files[9037] = "test_data_9037.txt";
test_data_files[9038] = "test_data_9038.txt";
test_data_files[9039] = "test_data_9039.txt";
test_data_files[9040] = "test_data_9040.txt";
test_data_files[9041] = "test_data_9041.txt";
test_data_files[9042] = "test_data_9042.txt";
test_data_files[9043] = "test_data_9043.txt";
test_data_files[9044] = "test_data_9044.txt";
test_data_files[9045] = "test_data_9045.txt";
test_data_files[9046] = "test_data_9046.txt";
test_data_files[9047] = "test_data_9047.txt";
test_data_files[9048] = "test_data_9048.txt";
test_data_files[9049] = "test_data_9049.txt";
test_data_files[9050] = "test_data_9050.txt";
test_data_files[9051] = "test_data_9051.txt";
test_data_files[9052] = "test_data_9052.txt";
test_data_files[9053] = "test_data_9053.txt";
test_data_files[9054] = "test_data_9054.txt";
test_data_files[9055] = "test_data_9055.txt";
test_data_files[9056] = "test_data_9056.txt";
test_data_files[9057] = "test_data_9057.txt";
test_data_files[9058] = "test_data_9058.txt";
test_data_files[9059] = "test_data_9059.txt";
test_data_files[9060] = "test_data_9060.txt";
test_data_files[9061] = "test_data_9061.txt";
test_data_files[9062] = "test_data_9062.txt";
test_data_files[9063] = "test_data_9063.txt";
test_data_files[9064] = "test_data_9064.txt";
test_data_files[9065] = "test_data_9065.txt";
test_data_files[9066] = "test_data_9066.txt";
test_data_files[9067] = "test_data_9067.txt";
test_data_files[9068] = "test_data_9068.txt";
test_data_files[9069] = "test_data_9069.txt";
test_data_files[9070] = "test_data_9070.txt";
test_data_files[9071] = "test_data_9071.txt";
test_data_files[9072] = "test_data_9072.txt";
test_data_files[9073] = "test_data_9073.txt";
test_data_files[9074] = "test_data_9074.txt";
test_data_files[9075] = "test_data_9075.txt";
test_data_files[9076] = "test_data_9076.txt";
test_data_files[9077] = "test_data_9077.txt";
test_data_files[9078] = "test_data_9078.txt";
test_data_files[9079] = "test_data_9079.txt";
test_data_files[9080] = "test_data_9080.txt";
test_data_files[9081] = "test_data_9081.txt";
test_data_files[9082] = "test_data_9082.txt";
test_data_files[9083] = "test_data_9083.txt";
test_data_files[9084] = "test_data_9084.txt";
test_data_files[9085] = "test_data_9085.txt";
test_data_files[9086] = "test_data_9086.txt";
test_data_files[9087] = "test_data_9087.txt";
test_data_files[9088] = "test_data_9088.txt";
test_data_files[9089] = "test_data_9089.txt";
test_data_files[9090] = "test_data_9090.txt";
test_data_files[9091] = "test_data_9091.txt";
test_data_files[9092] = "test_data_9092.txt";
test_data_files[9093] = "test_data_9093.txt";
test_data_files[9094] = "test_data_9094.txt";
test_data_files[9095] = "test_data_9095.txt";
test_data_files[9096] = "test_data_9096.txt";
test_data_files[9097] = "test_data_9097.txt";
test_data_files[9098] = "test_data_9098.txt";
test_data_files[9099] = "test_data_9099.txt";
test_data_files[9100] = "test_data_9100.txt";
test_data_files[9101] = "test_data_9101.txt";
test_data_files[9102] = "test_data_9102.txt";
test_data_files[9103] = "test_data_9103.txt";
test_data_files[9104] = "test_data_9104.txt";
test_data_files[9105] = "test_data_9105.txt";
test_data_files[9106] = "test_data_9106.txt";
test_data_files[9107] = "test_data_9107.txt";
test_data_files[9108] = "test_data_9108.txt";
test_data_files[9109] = "test_data_9109.txt";
test_data_files[9110] = "test_data_9110.txt";
test_data_files[9111] = "test_data_9111.txt";
test_data_files[9112] = "test_data_9112.txt";
test_data_files[9113] = "test_data_9113.txt";
test_data_files[9114] = "test_data_9114.txt";
test_data_files[9115] = "test_data_9115.txt";
test_data_files[9116] = "test_data_9116.txt";
test_data_files[9117] = "test_data_9117.txt";
test_data_files[9118] = "test_data_9118.txt";
test_data_files[9119] = "test_data_9119.txt";
test_data_files[9120] = "test_data_9120.txt";
test_data_files[9121] = "test_data_9121.txt";
test_data_files[9122] = "test_data_9122.txt";
test_data_files[9123] = "test_data_9123.txt";
test_data_files[9124] = "test_data_9124.txt";
test_data_files[9125] = "test_data_9125.txt";
test_data_files[9126] = "test_data_9126.txt";
test_data_files[9127] = "test_data_9127.txt";
test_data_files[9128] = "test_data_9128.txt";
test_data_files[9129] = "test_data_9129.txt";
test_data_files[9130] = "test_data_9130.txt";
test_data_files[9131] = "test_data_9131.txt";
test_data_files[9132] = "test_data_9132.txt";
test_data_files[9133] = "test_data_9133.txt";
test_data_files[9134] = "test_data_9134.txt";
test_data_files[9135] = "test_data_9135.txt";
test_data_files[9136] = "test_data_9136.txt";
test_data_files[9137] = "test_data_9137.txt";
test_data_files[9138] = "test_data_9138.txt";
test_data_files[9139] = "test_data_9139.txt";
test_data_files[9140] = "test_data_9140.txt";
test_data_files[9141] = "test_data_9141.txt";
test_data_files[9142] = "test_data_9142.txt";
test_data_files[9143] = "test_data_9143.txt";
test_data_files[9144] = "test_data_9144.txt";
test_data_files[9145] = "test_data_9145.txt";
test_data_files[9146] = "test_data_9146.txt";
test_data_files[9147] = "test_data_9147.txt";
test_data_files[9148] = "test_data_9148.txt";
test_data_files[9149] = "test_data_9149.txt";
test_data_files[9150] = "test_data_9150.txt";
test_data_files[9151] = "test_data_9151.txt";
test_data_files[9152] = "test_data_9152.txt";
test_data_files[9153] = "test_data_9153.txt";
test_data_files[9154] = "test_data_9154.txt";
test_data_files[9155] = "test_data_9155.txt";
test_data_files[9156] = "test_data_9156.txt";
test_data_files[9157] = "test_data_9157.txt";
test_data_files[9158] = "test_data_9158.txt";
test_data_files[9159] = "test_data_9159.txt";
test_data_files[9160] = "test_data_9160.txt";
test_data_files[9161] = "test_data_9161.txt";
test_data_files[9162] = "test_data_9162.txt";
test_data_files[9163] = "test_data_9163.txt";
test_data_files[9164] = "test_data_9164.txt";
test_data_files[9165] = "test_data_9165.txt";
test_data_files[9166] = "test_data_9166.txt";
test_data_files[9167] = "test_data_9167.txt";
test_data_files[9168] = "test_data_9168.txt";
test_data_files[9169] = "test_data_9169.txt";
test_data_files[9170] = "test_data_9170.txt";
test_data_files[9171] = "test_data_9171.txt";
test_data_files[9172] = "test_data_9172.txt";
test_data_files[9173] = "test_data_9173.txt";
test_data_files[9174] = "test_data_9174.txt";
test_data_files[9175] = "test_data_9175.txt";
test_data_files[9176] = "test_data_9176.txt";
test_data_files[9177] = "test_data_9177.txt";
test_data_files[9178] = "test_data_9178.txt";
test_data_files[9179] = "test_data_9179.txt";
test_data_files[9180] = "test_data_9180.txt";
test_data_files[9181] = "test_data_9181.txt";
test_data_files[9182] = "test_data_9182.txt";
test_data_files[9183] = "test_data_9183.txt";
test_data_files[9184] = "test_data_9184.txt";
test_data_files[9185] = "test_data_9185.txt";
test_data_files[9186] = "test_data_9186.txt";
test_data_files[9187] = "test_data_9187.txt";
test_data_files[9188] = "test_data_9188.txt";
test_data_files[9189] = "test_data_9189.txt";
test_data_files[9190] = "test_data_9190.txt";
test_data_files[9191] = "test_data_9191.txt";
test_data_files[9192] = "test_data_9192.txt";
test_data_files[9193] = "test_data_9193.txt";
test_data_files[9194] = "test_data_9194.txt";
test_data_files[9195] = "test_data_9195.txt";
test_data_files[9196] = "test_data_9196.txt";
test_data_files[9197] = "test_data_9197.txt";
test_data_files[9198] = "test_data_9198.txt";
test_data_files[9199] = "test_data_9199.txt";
test_data_files[9200] = "test_data_9200.txt";
test_data_files[9201] = "test_data_9201.txt";
test_data_files[9202] = "test_data_9202.txt";
test_data_files[9203] = "test_data_9203.txt";
test_data_files[9204] = "test_data_9204.txt";
test_data_files[9205] = "test_data_9205.txt";
test_data_files[9206] = "test_data_9206.txt";
test_data_files[9207] = "test_data_9207.txt";
test_data_files[9208] = "test_data_9208.txt";
test_data_files[9209] = "test_data_9209.txt";
test_data_files[9210] = "test_data_9210.txt";
test_data_files[9211] = "test_data_9211.txt";
test_data_files[9212] = "test_data_9212.txt";
test_data_files[9213] = "test_data_9213.txt";
test_data_files[9214] = "test_data_9214.txt";
test_data_files[9215] = "test_data_9215.txt";
test_data_files[9216] = "test_data_9216.txt";
test_data_files[9217] = "test_data_9217.txt";
test_data_files[9218] = "test_data_9218.txt";
test_data_files[9219] = "test_data_9219.txt";
test_data_files[9220] = "test_data_9220.txt";
test_data_files[9221] = "test_data_9221.txt";
test_data_files[9222] = "test_data_9222.txt";
test_data_files[9223] = "test_data_9223.txt";
test_data_files[9224] = "test_data_9224.txt";
test_data_files[9225] = "test_data_9225.txt";
test_data_files[9226] = "test_data_9226.txt";
test_data_files[9227] = "test_data_9227.txt";
test_data_files[9228] = "test_data_9228.txt";
test_data_files[9229] = "test_data_9229.txt";
test_data_files[9230] = "test_data_9230.txt";
test_data_files[9231] = "test_data_9231.txt";
test_data_files[9232] = "test_data_9232.txt";
test_data_files[9233] = "test_data_9233.txt";
test_data_files[9234] = "test_data_9234.txt";
test_data_files[9235] = "test_data_9235.txt";
test_data_files[9236] = "test_data_9236.txt";
test_data_files[9237] = "test_data_9237.txt";
test_data_files[9238] = "test_data_9238.txt";
test_data_files[9239] = "test_data_9239.txt";
test_data_files[9240] = "test_data_9240.txt";
test_data_files[9241] = "test_data_9241.txt";
test_data_files[9242] = "test_data_9242.txt";
test_data_files[9243] = "test_data_9243.txt";
test_data_files[9244] = "test_data_9244.txt";
test_data_files[9245] = "test_data_9245.txt";
test_data_files[9246] = "test_data_9246.txt";
test_data_files[9247] = "test_data_9247.txt";
test_data_files[9248] = "test_data_9248.txt";
test_data_files[9249] = "test_data_9249.txt";
test_data_files[9250] = "test_data_9250.txt";
test_data_files[9251] = "test_data_9251.txt";
test_data_files[9252] = "test_data_9252.txt";
test_data_files[9253] = "test_data_9253.txt";
test_data_files[9254] = "test_data_9254.txt";
test_data_files[9255] = "test_data_9255.txt";
test_data_files[9256] = "test_data_9256.txt";
test_data_files[9257] = "test_data_9257.txt";
test_data_files[9258] = "test_data_9258.txt";
test_data_files[9259] = "test_data_9259.txt";
test_data_files[9260] = "test_data_9260.txt";
test_data_files[9261] = "test_data_9261.txt";
test_data_files[9262] = "test_data_9262.txt";
test_data_files[9263] = "test_data_9263.txt";
test_data_files[9264] = "test_data_9264.txt";
test_data_files[9265] = "test_data_9265.txt";
test_data_files[9266] = "test_data_9266.txt";
test_data_files[9267] = "test_data_9267.txt";
test_data_files[9268] = "test_data_9268.txt";
test_data_files[9269] = "test_data_9269.txt";
test_data_files[9270] = "test_data_9270.txt";
test_data_files[9271] = "test_data_9271.txt";
test_data_files[9272] = "test_data_9272.txt";
test_data_files[9273] = "test_data_9273.txt";
test_data_files[9274] = "test_data_9274.txt";
test_data_files[9275] = "test_data_9275.txt";
test_data_files[9276] = "test_data_9276.txt";
test_data_files[9277] = "test_data_9277.txt";
test_data_files[9278] = "test_data_9278.txt";
test_data_files[9279] = "test_data_9279.txt";
test_data_files[9280] = "test_data_9280.txt";
test_data_files[9281] = "test_data_9281.txt";
test_data_files[9282] = "test_data_9282.txt";
test_data_files[9283] = "test_data_9283.txt";
test_data_files[9284] = "test_data_9284.txt";
test_data_files[9285] = "test_data_9285.txt";
test_data_files[9286] = "test_data_9286.txt";
test_data_files[9287] = "test_data_9287.txt";
test_data_files[9288] = "test_data_9288.txt";
test_data_files[9289] = "test_data_9289.txt";
test_data_files[9290] = "test_data_9290.txt";
test_data_files[9291] = "test_data_9291.txt";
test_data_files[9292] = "test_data_9292.txt";
test_data_files[9293] = "test_data_9293.txt";
test_data_files[9294] = "test_data_9294.txt";
test_data_files[9295] = "test_data_9295.txt";
test_data_files[9296] = "test_data_9296.txt";
test_data_files[9297] = "test_data_9297.txt";
test_data_files[9298] = "test_data_9298.txt";
test_data_files[9299] = "test_data_9299.txt";
test_data_files[9300] = "test_data_9300.txt";
test_data_files[9301] = "test_data_9301.txt";
test_data_files[9302] = "test_data_9302.txt";
test_data_files[9303] = "test_data_9303.txt";
test_data_files[9304] = "test_data_9304.txt";
test_data_files[9305] = "test_data_9305.txt";
test_data_files[9306] = "test_data_9306.txt";
test_data_files[9307] = "test_data_9307.txt";
test_data_files[9308] = "test_data_9308.txt";
test_data_files[9309] = "test_data_9309.txt";
test_data_files[9310] = "test_data_9310.txt";
test_data_files[9311] = "test_data_9311.txt";
test_data_files[9312] = "test_data_9312.txt";
test_data_files[9313] = "test_data_9313.txt";
test_data_files[9314] = "test_data_9314.txt";
test_data_files[9315] = "test_data_9315.txt";
test_data_files[9316] = "test_data_9316.txt";
test_data_files[9317] = "test_data_9317.txt";
test_data_files[9318] = "test_data_9318.txt";
test_data_files[9319] = "test_data_9319.txt";
test_data_files[9320] = "test_data_9320.txt";
test_data_files[9321] = "test_data_9321.txt";
test_data_files[9322] = "test_data_9322.txt";
test_data_files[9323] = "test_data_9323.txt";
test_data_files[9324] = "test_data_9324.txt";
test_data_files[9325] = "test_data_9325.txt";
test_data_files[9326] = "test_data_9326.txt";
test_data_files[9327] = "test_data_9327.txt";
test_data_files[9328] = "test_data_9328.txt";
test_data_files[9329] = "test_data_9329.txt";
test_data_files[9330] = "test_data_9330.txt";
test_data_files[9331] = "test_data_9331.txt";
test_data_files[9332] = "test_data_9332.txt";
test_data_files[9333] = "test_data_9333.txt";
test_data_files[9334] = "test_data_9334.txt";
test_data_files[9335] = "test_data_9335.txt";
test_data_files[9336] = "test_data_9336.txt";
test_data_files[9337] = "test_data_9337.txt";
test_data_files[9338] = "test_data_9338.txt";
test_data_files[9339] = "test_data_9339.txt";
test_data_files[9340] = "test_data_9340.txt";
test_data_files[9341] = "test_data_9341.txt";
test_data_files[9342] = "test_data_9342.txt";
test_data_files[9343] = "test_data_9343.txt";
test_data_files[9344] = "test_data_9344.txt";
test_data_files[9345] = "test_data_9345.txt";
test_data_files[9346] = "test_data_9346.txt";
test_data_files[9347] = "test_data_9347.txt";
test_data_files[9348] = "test_data_9348.txt";
test_data_files[9349] = "test_data_9349.txt";
test_data_files[9350] = "test_data_9350.txt";
test_data_files[9351] = "test_data_9351.txt";
test_data_files[9352] = "test_data_9352.txt";
test_data_files[9353] = "test_data_9353.txt";
test_data_files[9354] = "test_data_9354.txt";
test_data_files[9355] = "test_data_9355.txt";
test_data_files[9356] = "test_data_9356.txt";
test_data_files[9357] = "test_data_9357.txt";
test_data_files[9358] = "test_data_9358.txt";
test_data_files[9359] = "test_data_9359.txt";
test_data_files[9360] = "test_data_9360.txt";
test_data_files[9361] = "test_data_9361.txt";
test_data_files[9362] = "test_data_9362.txt";
test_data_files[9363] = "test_data_9363.txt";
test_data_files[9364] = "test_data_9364.txt";
test_data_files[9365] = "test_data_9365.txt";
test_data_files[9366] = "test_data_9366.txt";
test_data_files[9367] = "test_data_9367.txt";
test_data_files[9368] = "test_data_9368.txt";
test_data_files[9369] = "test_data_9369.txt";
test_data_files[9370] = "test_data_9370.txt";
test_data_files[9371] = "test_data_9371.txt";
test_data_files[9372] = "test_data_9372.txt";
test_data_files[9373] = "test_data_9373.txt";
test_data_files[9374] = "test_data_9374.txt";
test_data_files[9375] = "test_data_9375.txt";
test_data_files[9376] = "test_data_9376.txt";
test_data_files[9377] = "test_data_9377.txt";
test_data_files[9378] = "test_data_9378.txt";
test_data_files[9379] = "test_data_9379.txt";
test_data_files[9380] = "test_data_9380.txt";
test_data_files[9381] = "test_data_9381.txt";
test_data_files[9382] = "test_data_9382.txt";
test_data_files[9383] = "test_data_9383.txt";
test_data_files[9384] = "test_data_9384.txt";
test_data_files[9385] = "test_data_9385.txt";
test_data_files[9386] = "test_data_9386.txt";
test_data_files[9387] = "test_data_9387.txt";
test_data_files[9388] = "test_data_9388.txt";
test_data_files[9389] = "test_data_9389.txt";
test_data_files[9390] = "test_data_9390.txt";
test_data_files[9391] = "test_data_9391.txt";
test_data_files[9392] = "test_data_9392.txt";
test_data_files[9393] = "test_data_9393.txt";
test_data_files[9394] = "test_data_9394.txt";
test_data_files[9395] = "test_data_9395.txt";
test_data_files[9396] = "test_data_9396.txt";
test_data_files[9397] = "test_data_9397.txt";
test_data_files[9398] = "test_data_9398.txt";
test_data_files[9399] = "test_data_9399.txt";
test_data_files[9400] = "test_data_9400.txt";
test_data_files[9401] = "test_data_9401.txt";
test_data_files[9402] = "test_data_9402.txt";
test_data_files[9403] = "test_data_9403.txt";
test_data_files[9404] = "test_data_9404.txt";
test_data_files[9405] = "test_data_9405.txt";
test_data_files[9406] = "test_data_9406.txt";
test_data_files[9407] = "test_data_9407.txt";
test_data_files[9408] = "test_data_9408.txt";
test_data_files[9409] = "test_data_9409.txt";
test_data_files[9410] = "test_data_9410.txt";
test_data_files[9411] = "test_data_9411.txt";
test_data_files[9412] = "test_data_9412.txt";
test_data_files[9413] = "test_data_9413.txt";
test_data_files[9414] = "test_data_9414.txt";
test_data_files[9415] = "test_data_9415.txt";
test_data_files[9416] = "test_data_9416.txt";
test_data_files[9417] = "test_data_9417.txt";
test_data_files[9418] = "test_data_9418.txt";
test_data_files[9419] = "test_data_9419.txt";
test_data_files[9420] = "test_data_9420.txt";
test_data_files[9421] = "test_data_9421.txt";
test_data_files[9422] = "test_data_9422.txt";
test_data_files[9423] = "test_data_9423.txt";
test_data_files[9424] = "test_data_9424.txt";
test_data_files[9425] = "test_data_9425.txt";
test_data_files[9426] = "test_data_9426.txt";
test_data_files[9427] = "test_data_9427.txt";
test_data_files[9428] = "test_data_9428.txt";
test_data_files[9429] = "test_data_9429.txt";
test_data_files[9430] = "test_data_9430.txt";
test_data_files[9431] = "test_data_9431.txt";
test_data_files[9432] = "test_data_9432.txt";
test_data_files[9433] = "test_data_9433.txt";
test_data_files[9434] = "test_data_9434.txt";
test_data_files[9435] = "test_data_9435.txt";
test_data_files[9436] = "test_data_9436.txt";
test_data_files[9437] = "test_data_9437.txt";
test_data_files[9438] = "test_data_9438.txt";
test_data_files[9439] = "test_data_9439.txt";
test_data_files[9440] = "test_data_9440.txt";
test_data_files[9441] = "test_data_9441.txt";
test_data_files[9442] = "test_data_9442.txt";
test_data_files[9443] = "test_data_9443.txt";
test_data_files[9444] = "test_data_9444.txt";
test_data_files[9445] = "test_data_9445.txt";
test_data_files[9446] = "test_data_9446.txt";
test_data_files[9447] = "test_data_9447.txt";
test_data_files[9448] = "test_data_9448.txt";
test_data_files[9449] = "test_data_9449.txt";
test_data_files[9450] = "test_data_9450.txt";
test_data_files[9451] = "test_data_9451.txt";
test_data_files[9452] = "test_data_9452.txt";
test_data_files[9453] = "test_data_9453.txt";
test_data_files[9454] = "test_data_9454.txt";
test_data_files[9455] = "test_data_9455.txt";
test_data_files[9456] = "test_data_9456.txt";
test_data_files[9457] = "test_data_9457.txt";
test_data_files[9458] = "test_data_9458.txt";
test_data_files[9459] = "test_data_9459.txt";
test_data_files[9460] = "test_data_9460.txt";
test_data_files[9461] = "test_data_9461.txt";
test_data_files[9462] = "test_data_9462.txt";
test_data_files[9463] = "test_data_9463.txt";
test_data_files[9464] = "test_data_9464.txt";
test_data_files[9465] = "test_data_9465.txt";
test_data_files[9466] = "test_data_9466.txt";
test_data_files[9467] = "test_data_9467.txt";
test_data_files[9468] = "test_data_9468.txt";
test_data_files[9469] = "test_data_9469.txt";
test_data_files[9470] = "test_data_9470.txt";
test_data_files[9471] = "test_data_9471.txt";
test_data_files[9472] = "test_data_9472.txt";
test_data_files[9473] = "test_data_9473.txt";
test_data_files[9474] = "test_data_9474.txt";
test_data_files[9475] = "test_data_9475.txt";
test_data_files[9476] = "test_data_9476.txt";
test_data_files[9477] = "test_data_9477.txt";
test_data_files[9478] = "test_data_9478.txt";
test_data_files[9479] = "test_data_9479.txt";
test_data_files[9480] = "test_data_9480.txt";
test_data_files[9481] = "test_data_9481.txt";
test_data_files[9482] = "test_data_9482.txt";
test_data_files[9483] = "test_data_9483.txt";
test_data_files[9484] = "test_data_9484.txt";
test_data_files[9485] = "test_data_9485.txt";
test_data_files[9486] = "test_data_9486.txt";
test_data_files[9487] = "test_data_9487.txt";
test_data_files[9488] = "test_data_9488.txt";
test_data_files[9489] = "test_data_9489.txt";
test_data_files[9490] = "test_data_9490.txt";
test_data_files[9491] = "test_data_9491.txt";
test_data_files[9492] = "test_data_9492.txt";
test_data_files[9493] = "test_data_9493.txt";
test_data_files[9494] = "test_data_9494.txt";
test_data_files[9495] = "test_data_9495.txt";
test_data_files[9496] = "test_data_9496.txt";
test_data_files[9497] = "test_data_9497.txt";
test_data_files[9498] = "test_data_9498.txt";
test_data_files[9499] = "test_data_9499.txt";
test_data_files[9500] = "test_data_9500.txt";
test_data_files[9501] = "test_data_9501.txt";
test_data_files[9502] = "test_data_9502.txt";
test_data_files[9503] = "test_data_9503.txt";
test_data_files[9504] = "test_data_9504.txt";
test_data_files[9505] = "test_data_9505.txt";
test_data_files[9506] = "test_data_9506.txt";
test_data_files[9507] = "test_data_9507.txt";
test_data_files[9508] = "test_data_9508.txt";
test_data_files[9509] = "test_data_9509.txt";
test_data_files[9510] = "test_data_9510.txt";
test_data_files[9511] = "test_data_9511.txt";
test_data_files[9512] = "test_data_9512.txt";
test_data_files[9513] = "test_data_9513.txt";
test_data_files[9514] = "test_data_9514.txt";
test_data_files[9515] = "test_data_9515.txt";
test_data_files[9516] = "test_data_9516.txt";
test_data_files[9517] = "test_data_9517.txt";
test_data_files[9518] = "test_data_9518.txt";
test_data_files[9519] = "test_data_9519.txt";
test_data_files[9520] = "test_data_9520.txt";
test_data_files[9521] = "test_data_9521.txt";
test_data_files[9522] = "test_data_9522.txt";
test_data_files[9523] = "test_data_9523.txt";
test_data_files[9524] = "test_data_9524.txt";
test_data_files[9525] = "test_data_9525.txt";
test_data_files[9526] = "test_data_9526.txt";
test_data_files[9527] = "test_data_9527.txt";
test_data_files[9528] = "test_data_9528.txt";
test_data_files[9529] = "test_data_9529.txt";
test_data_files[9530] = "test_data_9530.txt";
test_data_files[9531] = "test_data_9531.txt";
test_data_files[9532] = "test_data_9532.txt";
test_data_files[9533] = "test_data_9533.txt";
test_data_files[9534] = "test_data_9534.txt";
test_data_files[9535] = "test_data_9535.txt";
test_data_files[9536] = "test_data_9536.txt";
test_data_files[9537] = "test_data_9537.txt";
test_data_files[9538] = "test_data_9538.txt";
test_data_files[9539] = "test_data_9539.txt";
test_data_files[9540] = "test_data_9540.txt";
test_data_files[9541] = "test_data_9541.txt";
test_data_files[9542] = "test_data_9542.txt";
test_data_files[9543] = "test_data_9543.txt";
test_data_files[9544] = "test_data_9544.txt";
test_data_files[9545] = "test_data_9545.txt";
test_data_files[9546] = "test_data_9546.txt";
test_data_files[9547] = "test_data_9547.txt";
test_data_files[9548] = "test_data_9548.txt";
test_data_files[9549] = "test_data_9549.txt";
test_data_files[9550] = "test_data_9550.txt";
test_data_files[9551] = "test_data_9551.txt";
test_data_files[9552] = "test_data_9552.txt";
test_data_files[9553] = "test_data_9553.txt";
test_data_files[9554] = "test_data_9554.txt";
test_data_files[9555] = "test_data_9555.txt";
test_data_files[9556] = "test_data_9556.txt";
test_data_files[9557] = "test_data_9557.txt";
test_data_files[9558] = "test_data_9558.txt";
test_data_files[9559] = "test_data_9559.txt";
test_data_files[9560] = "test_data_9560.txt";
test_data_files[9561] = "test_data_9561.txt";
test_data_files[9562] = "test_data_9562.txt";
test_data_files[9563] = "test_data_9563.txt";
test_data_files[9564] = "test_data_9564.txt";
test_data_files[9565] = "test_data_9565.txt";
test_data_files[9566] = "test_data_9566.txt";
test_data_files[9567] = "test_data_9567.txt";
test_data_files[9568] = "test_data_9568.txt";
test_data_files[9569] = "test_data_9569.txt";
test_data_files[9570] = "test_data_9570.txt";
test_data_files[9571] = "test_data_9571.txt";
test_data_files[9572] = "test_data_9572.txt";
test_data_files[9573] = "test_data_9573.txt";
test_data_files[9574] = "test_data_9574.txt";
test_data_files[9575] = "test_data_9575.txt";
test_data_files[9576] = "test_data_9576.txt";
test_data_files[9577] = "test_data_9577.txt";
test_data_files[9578] = "test_data_9578.txt";
test_data_files[9579] = "test_data_9579.txt";
test_data_files[9580] = "test_data_9580.txt";
test_data_files[9581] = "test_data_9581.txt";
test_data_files[9582] = "test_data_9582.txt";
test_data_files[9583] = "test_data_9583.txt";
test_data_files[9584] = "test_data_9584.txt";
test_data_files[9585] = "test_data_9585.txt";
test_data_files[9586] = "test_data_9586.txt";
test_data_files[9587] = "test_data_9587.txt";
test_data_files[9588] = "test_data_9588.txt";
test_data_files[9589] = "test_data_9589.txt";
test_data_files[9590] = "test_data_9590.txt";
test_data_files[9591] = "test_data_9591.txt";
test_data_files[9592] = "test_data_9592.txt";
test_data_files[9593] = "test_data_9593.txt";
test_data_files[9594] = "test_data_9594.txt";
test_data_files[9595] = "test_data_9595.txt";
test_data_files[9596] = "test_data_9596.txt";
test_data_files[9597] = "test_data_9597.txt";
test_data_files[9598] = "test_data_9598.txt";
test_data_files[9599] = "test_data_9599.txt";
test_data_files[9600] = "test_data_9600.txt";
test_data_files[9601] = "test_data_9601.txt";
test_data_files[9602] = "test_data_9602.txt";
test_data_files[9603] = "test_data_9603.txt";
test_data_files[9604] = "test_data_9604.txt";
test_data_files[9605] = "test_data_9605.txt";
test_data_files[9606] = "test_data_9606.txt";
test_data_files[9607] = "test_data_9607.txt";
test_data_files[9608] = "test_data_9608.txt";
test_data_files[9609] = "test_data_9609.txt";
test_data_files[9610] = "test_data_9610.txt";
test_data_files[9611] = "test_data_9611.txt";
test_data_files[9612] = "test_data_9612.txt";
test_data_files[9613] = "test_data_9613.txt";
test_data_files[9614] = "test_data_9614.txt";
test_data_files[9615] = "test_data_9615.txt";
test_data_files[9616] = "test_data_9616.txt";
test_data_files[9617] = "test_data_9617.txt";
test_data_files[9618] = "test_data_9618.txt";
test_data_files[9619] = "test_data_9619.txt";
test_data_files[9620] = "test_data_9620.txt";
test_data_files[9621] = "test_data_9621.txt";
test_data_files[9622] = "test_data_9622.txt";
test_data_files[9623] = "test_data_9623.txt";
test_data_files[9624] = "test_data_9624.txt";
test_data_files[9625] = "test_data_9625.txt";
test_data_files[9626] = "test_data_9626.txt";
test_data_files[9627] = "test_data_9627.txt";
test_data_files[9628] = "test_data_9628.txt";
test_data_files[9629] = "test_data_9629.txt";
test_data_files[9630] = "test_data_9630.txt";
test_data_files[9631] = "test_data_9631.txt";
test_data_files[9632] = "test_data_9632.txt";
test_data_files[9633] = "test_data_9633.txt";
test_data_files[9634] = "test_data_9634.txt";
test_data_files[9635] = "test_data_9635.txt";
test_data_files[9636] = "test_data_9636.txt";
test_data_files[9637] = "test_data_9637.txt";
test_data_files[9638] = "test_data_9638.txt";
test_data_files[9639] = "test_data_9639.txt";
test_data_files[9640] = "test_data_9640.txt";
test_data_files[9641] = "test_data_9641.txt";
test_data_files[9642] = "test_data_9642.txt";
test_data_files[9643] = "test_data_9643.txt";
test_data_files[9644] = "test_data_9644.txt";
test_data_files[9645] = "test_data_9645.txt";
test_data_files[9646] = "test_data_9646.txt";
test_data_files[9647] = "test_data_9647.txt";
test_data_files[9648] = "test_data_9648.txt";
test_data_files[9649] = "test_data_9649.txt";
test_data_files[9650] = "test_data_9650.txt";
test_data_files[9651] = "test_data_9651.txt";
test_data_files[9652] = "test_data_9652.txt";
test_data_files[9653] = "test_data_9653.txt";
test_data_files[9654] = "test_data_9654.txt";
test_data_files[9655] = "test_data_9655.txt";
test_data_files[9656] = "test_data_9656.txt";
test_data_files[9657] = "test_data_9657.txt";
test_data_files[9658] = "test_data_9658.txt";
test_data_files[9659] = "test_data_9659.txt";
test_data_files[9660] = "test_data_9660.txt";
test_data_files[9661] = "test_data_9661.txt";
test_data_files[9662] = "test_data_9662.txt";
test_data_files[9663] = "test_data_9663.txt";
test_data_files[9664] = "test_data_9664.txt";
test_data_files[9665] = "test_data_9665.txt";
test_data_files[9666] = "test_data_9666.txt";
test_data_files[9667] = "test_data_9667.txt";
test_data_files[9668] = "test_data_9668.txt";
test_data_files[9669] = "test_data_9669.txt";
test_data_files[9670] = "test_data_9670.txt";
test_data_files[9671] = "test_data_9671.txt";
test_data_files[9672] = "test_data_9672.txt";
test_data_files[9673] = "test_data_9673.txt";
test_data_files[9674] = "test_data_9674.txt";
test_data_files[9675] = "test_data_9675.txt";
test_data_files[9676] = "test_data_9676.txt";
test_data_files[9677] = "test_data_9677.txt";
test_data_files[9678] = "test_data_9678.txt";
test_data_files[9679] = "test_data_9679.txt";
test_data_files[9680] = "test_data_9680.txt";
test_data_files[9681] = "test_data_9681.txt";
test_data_files[9682] = "test_data_9682.txt";
test_data_files[9683] = "test_data_9683.txt";
test_data_files[9684] = "test_data_9684.txt";
test_data_files[9685] = "test_data_9685.txt";
test_data_files[9686] = "test_data_9686.txt";
test_data_files[9687] = "test_data_9687.txt";
test_data_files[9688] = "test_data_9688.txt";
test_data_files[9689] = "test_data_9689.txt";
test_data_files[9690] = "test_data_9690.txt";
test_data_files[9691] = "test_data_9691.txt";
test_data_files[9692] = "test_data_9692.txt";
test_data_files[9693] = "test_data_9693.txt";
test_data_files[9694] = "test_data_9694.txt";
test_data_files[9695] = "test_data_9695.txt";
test_data_files[9696] = "test_data_9696.txt";
test_data_files[9697] = "test_data_9697.txt";
test_data_files[9698] = "test_data_9698.txt";
test_data_files[9699] = "test_data_9699.txt";
test_data_files[9700] = "test_data_9700.txt";
test_data_files[9701] = "test_data_9701.txt";
test_data_files[9702] = "test_data_9702.txt";
test_data_files[9703] = "test_data_9703.txt";
test_data_files[9704] = "test_data_9704.txt";
test_data_files[9705] = "test_data_9705.txt";
test_data_files[9706] = "test_data_9706.txt";
test_data_files[9707] = "test_data_9707.txt";
test_data_files[9708] = "test_data_9708.txt";
test_data_files[9709] = "test_data_9709.txt";
test_data_files[9710] = "test_data_9710.txt";
test_data_files[9711] = "test_data_9711.txt";
test_data_files[9712] = "test_data_9712.txt";
test_data_files[9713] = "test_data_9713.txt";
test_data_files[9714] = "test_data_9714.txt";
test_data_files[9715] = "test_data_9715.txt";
test_data_files[9716] = "test_data_9716.txt";
test_data_files[9717] = "test_data_9717.txt";
test_data_files[9718] = "test_data_9718.txt";
test_data_files[9719] = "test_data_9719.txt";
test_data_files[9720] = "test_data_9720.txt";
test_data_files[9721] = "test_data_9721.txt";
test_data_files[9722] = "test_data_9722.txt";
test_data_files[9723] = "test_data_9723.txt";
test_data_files[9724] = "test_data_9724.txt";
test_data_files[9725] = "test_data_9725.txt";
test_data_files[9726] = "test_data_9726.txt";
test_data_files[9727] = "test_data_9727.txt";
test_data_files[9728] = "test_data_9728.txt";
test_data_files[9729] = "test_data_9729.txt";
test_data_files[9730] = "test_data_9730.txt";
test_data_files[9731] = "test_data_9731.txt";
test_data_files[9732] = "test_data_9732.txt";
test_data_files[9733] = "test_data_9733.txt";
test_data_files[9734] = "test_data_9734.txt";
test_data_files[9735] = "test_data_9735.txt";
test_data_files[9736] = "test_data_9736.txt";
test_data_files[9737] = "test_data_9737.txt";
test_data_files[9738] = "test_data_9738.txt";
test_data_files[9739] = "test_data_9739.txt";
test_data_files[9740] = "test_data_9740.txt";
test_data_files[9741] = "test_data_9741.txt";
test_data_files[9742] = "test_data_9742.txt";
test_data_files[9743] = "test_data_9743.txt";
test_data_files[9744] = "test_data_9744.txt";
test_data_files[9745] = "test_data_9745.txt";
test_data_files[9746] = "test_data_9746.txt";
test_data_files[9747] = "test_data_9747.txt";
test_data_files[9748] = "test_data_9748.txt";
test_data_files[9749] = "test_data_9749.txt";
test_data_files[9750] = "test_data_9750.txt";
test_data_files[9751] = "test_data_9751.txt";
test_data_files[9752] = "test_data_9752.txt";
test_data_files[9753] = "test_data_9753.txt";
test_data_files[9754] = "test_data_9754.txt";
test_data_files[9755] = "test_data_9755.txt";
test_data_files[9756] = "test_data_9756.txt";
test_data_files[9757] = "test_data_9757.txt";
test_data_files[9758] = "test_data_9758.txt";
test_data_files[9759] = "test_data_9759.txt";
test_data_files[9760] = "test_data_9760.txt";
test_data_files[9761] = "test_data_9761.txt";
test_data_files[9762] = "test_data_9762.txt";
test_data_files[9763] = "test_data_9763.txt";
test_data_files[9764] = "test_data_9764.txt";
test_data_files[9765] = "test_data_9765.txt";
test_data_files[9766] = "test_data_9766.txt";
test_data_files[9767] = "test_data_9767.txt";
test_data_files[9768] = "test_data_9768.txt";
test_data_files[9769] = "test_data_9769.txt";
test_data_files[9770] = "test_data_9770.txt";
test_data_files[9771] = "test_data_9771.txt";
test_data_files[9772] = "test_data_9772.txt";
test_data_files[9773] = "test_data_9773.txt";
test_data_files[9774] = "test_data_9774.txt";
test_data_files[9775] = "test_data_9775.txt";
test_data_files[9776] = "test_data_9776.txt";
test_data_files[9777] = "test_data_9777.txt";
test_data_files[9778] = "test_data_9778.txt";
test_data_files[9779] = "test_data_9779.txt";
test_data_files[9780] = "test_data_9780.txt";
test_data_files[9781] = "test_data_9781.txt";
test_data_files[9782] = "test_data_9782.txt";
test_data_files[9783] = "test_data_9783.txt";
test_data_files[9784] = "test_data_9784.txt";
test_data_files[9785] = "test_data_9785.txt";
test_data_files[9786] = "test_data_9786.txt";
test_data_files[9787] = "test_data_9787.txt";
test_data_files[9788] = "test_data_9788.txt";
test_data_files[9789] = "test_data_9789.txt";
test_data_files[9790] = "test_data_9790.txt";
test_data_files[9791] = "test_data_9791.txt";
test_data_files[9792] = "test_data_9792.txt";
test_data_files[9793] = "test_data_9793.txt";
test_data_files[9794] = "test_data_9794.txt";
test_data_files[9795] = "test_data_9795.txt";
test_data_files[9796] = "test_data_9796.txt";
test_data_files[9797] = "test_data_9797.txt";
test_data_files[9798] = "test_data_9798.txt";
test_data_files[9799] = "test_data_9799.txt";
test_data_files[9800] = "test_data_9800.txt";
test_data_files[9801] = "test_data_9801.txt";
test_data_files[9802] = "test_data_9802.txt";
test_data_files[9803] = "test_data_9803.txt";
test_data_files[9804] = "test_data_9804.txt";
test_data_files[9805] = "test_data_9805.txt";
test_data_files[9806] = "test_data_9806.txt";
test_data_files[9807] = "test_data_9807.txt";
test_data_files[9808] = "test_data_9808.txt";
test_data_files[9809] = "test_data_9809.txt";
test_data_files[9810] = "test_data_9810.txt";
test_data_files[9811] = "test_data_9811.txt";
test_data_files[9812] = "test_data_9812.txt";
test_data_files[9813] = "test_data_9813.txt";
test_data_files[9814] = "test_data_9814.txt";
test_data_files[9815] = "test_data_9815.txt";
test_data_files[9816] = "test_data_9816.txt";
test_data_files[9817] = "test_data_9817.txt";
test_data_files[9818] = "test_data_9818.txt";
test_data_files[9819] = "test_data_9819.txt";
test_data_files[9820] = "test_data_9820.txt";
test_data_files[9821] = "test_data_9821.txt";
test_data_files[9822] = "test_data_9822.txt";
test_data_files[9823] = "test_data_9823.txt";
test_data_files[9824] = "test_data_9824.txt";
test_data_files[9825] = "test_data_9825.txt";
test_data_files[9826] = "test_data_9826.txt";
test_data_files[9827] = "test_data_9827.txt";
test_data_files[9828] = "test_data_9828.txt";
test_data_files[9829] = "test_data_9829.txt";
test_data_files[9830] = "test_data_9830.txt";
test_data_files[9831] = "test_data_9831.txt";
test_data_files[9832] = "test_data_9832.txt";
test_data_files[9833] = "test_data_9833.txt";
test_data_files[9834] = "test_data_9834.txt";
test_data_files[9835] = "test_data_9835.txt";
test_data_files[9836] = "test_data_9836.txt";
test_data_files[9837] = "test_data_9837.txt";
test_data_files[9838] = "test_data_9838.txt";
test_data_files[9839] = "test_data_9839.txt";
test_data_files[9840] = "test_data_9840.txt";
test_data_files[9841] = "test_data_9841.txt";
test_data_files[9842] = "test_data_9842.txt";
test_data_files[9843] = "test_data_9843.txt";
test_data_files[9844] = "test_data_9844.txt";
test_data_files[9845] = "test_data_9845.txt";
test_data_files[9846] = "test_data_9846.txt";
test_data_files[9847] = "test_data_9847.txt";
test_data_files[9848] = "test_data_9848.txt";
test_data_files[9849] = "test_data_9849.txt";
test_data_files[9850] = "test_data_9850.txt";
test_data_files[9851] = "test_data_9851.txt";
test_data_files[9852] = "test_data_9852.txt";
test_data_files[9853] = "test_data_9853.txt";
test_data_files[9854] = "test_data_9854.txt";
test_data_files[9855] = "test_data_9855.txt";
test_data_files[9856] = "test_data_9856.txt";
test_data_files[9857] = "test_data_9857.txt";
test_data_files[9858] = "test_data_9858.txt";
test_data_files[9859] = "test_data_9859.txt";
test_data_files[9860] = "test_data_9860.txt";
test_data_files[9861] = "test_data_9861.txt";
test_data_files[9862] = "test_data_9862.txt";
test_data_files[9863] = "test_data_9863.txt";
test_data_files[9864] = "test_data_9864.txt";
test_data_files[9865] = "test_data_9865.txt";
test_data_files[9866] = "test_data_9866.txt";
test_data_files[9867] = "test_data_9867.txt";
test_data_files[9868] = "test_data_9868.txt";
test_data_files[9869] = "test_data_9869.txt";
test_data_files[9870] = "test_data_9870.txt";
test_data_files[9871] = "test_data_9871.txt";
test_data_files[9872] = "test_data_9872.txt";
test_data_files[9873] = "test_data_9873.txt";
test_data_files[9874] = "test_data_9874.txt";
test_data_files[9875] = "test_data_9875.txt";
test_data_files[9876] = "test_data_9876.txt";
test_data_files[9877] = "test_data_9877.txt";
test_data_files[9878] = "test_data_9878.txt";
test_data_files[9879] = "test_data_9879.txt";
test_data_files[9880] = "test_data_9880.txt";
test_data_files[9881] = "test_data_9881.txt";
test_data_files[9882] = "test_data_9882.txt";
test_data_files[9883] = "test_data_9883.txt";
test_data_files[9884] = "test_data_9884.txt";
test_data_files[9885] = "test_data_9885.txt";
test_data_files[9886] = "test_data_9886.txt";
test_data_files[9887] = "test_data_9887.txt";
test_data_files[9888] = "test_data_9888.txt";
test_data_files[9889] = "test_data_9889.txt";
test_data_files[9890] = "test_data_9890.txt";
test_data_files[9891] = "test_data_9891.txt";
test_data_files[9892] = "test_data_9892.txt";
test_data_files[9893] = "test_data_9893.txt";
test_data_files[9894] = "test_data_9894.txt";
test_data_files[9895] = "test_data_9895.txt";
test_data_files[9896] = "test_data_9896.txt";
test_data_files[9897] = "test_data_9897.txt";
test_data_files[9898] = "test_data_9898.txt";
test_data_files[9899] = "test_data_9899.txt";
test_data_files[9900] = "test_data_9900.txt";
test_data_files[9901] = "test_data_9901.txt";
test_data_files[9902] = "test_data_9902.txt";
test_data_files[9903] = "test_data_9903.txt";
test_data_files[9904] = "test_data_9904.txt";
test_data_files[9905] = "test_data_9905.txt";
test_data_files[9906] = "test_data_9906.txt";
test_data_files[9907] = "test_data_9907.txt";
test_data_files[9908] = "test_data_9908.txt";
test_data_files[9909] = "test_data_9909.txt";
test_data_files[9910] = "test_data_9910.txt";
test_data_files[9911] = "test_data_9911.txt";
test_data_files[9912] = "test_data_9912.txt";
test_data_files[9913] = "test_data_9913.txt";
test_data_files[9914] = "test_data_9914.txt";
test_data_files[9915] = "test_data_9915.txt";
test_data_files[9916] = "test_data_9916.txt";
test_data_files[9917] = "test_data_9917.txt";
test_data_files[9918] = "test_data_9918.txt";
test_data_files[9919] = "test_data_9919.txt";
test_data_files[9920] = "test_data_9920.txt";
test_data_files[9921] = "test_data_9921.txt";
test_data_files[9922] = "test_data_9922.txt";
test_data_files[9923] = "test_data_9923.txt";
test_data_files[9924] = "test_data_9924.txt";
test_data_files[9925] = "test_data_9925.txt";
test_data_files[9926] = "test_data_9926.txt";
test_data_files[9927] = "test_data_9927.txt";
test_data_files[9928] = "test_data_9928.txt";
test_data_files[9929] = "test_data_9929.txt";
test_data_files[9930] = "test_data_9930.txt";
test_data_files[9931] = "test_data_9931.txt";
test_data_files[9932] = "test_data_9932.txt";
test_data_files[9933] = "test_data_9933.txt";
test_data_files[9934] = "test_data_9934.txt";
test_data_files[9935] = "test_data_9935.txt";
test_data_files[9936] = "test_data_9936.txt";
test_data_files[9937] = "test_data_9937.txt";
test_data_files[9938] = "test_data_9938.txt";
test_data_files[9939] = "test_data_9939.txt";
test_data_files[9940] = "test_data_9940.txt";
test_data_files[9941] = "test_data_9941.txt";
test_data_files[9942] = "test_data_9942.txt";
test_data_files[9943] = "test_data_9943.txt";
test_data_files[9944] = "test_data_9944.txt";
test_data_files[9945] = "test_data_9945.txt";
test_data_files[9946] = "test_data_9946.txt";
test_data_files[9947] = "test_data_9947.txt";
test_data_files[9948] = "test_data_9948.txt";
test_data_files[9949] = "test_data_9949.txt";
test_data_files[9950] = "test_data_9950.txt";
test_data_files[9951] = "test_data_9951.txt";
test_data_files[9952] = "test_data_9952.txt";
test_data_files[9953] = "test_data_9953.txt";
test_data_files[9954] = "test_data_9954.txt";
test_data_files[9955] = "test_data_9955.txt";
test_data_files[9956] = "test_data_9956.txt";
test_data_files[9957] = "test_data_9957.txt";
test_data_files[9958] = "test_data_9958.txt";
test_data_files[9959] = "test_data_9959.txt";
test_data_files[9960] = "test_data_9960.txt";
test_data_files[9961] = "test_data_9961.txt";
test_data_files[9962] = "test_data_9962.txt";
test_data_files[9963] = "test_data_9963.txt";
test_data_files[9964] = "test_data_9964.txt";
test_data_files[9965] = "test_data_9965.txt";
test_data_files[9966] = "test_data_9966.txt";
test_data_files[9967] = "test_data_9967.txt";
test_data_files[9968] = "test_data_9968.txt";
test_data_files[9969] = "test_data_9969.txt";
test_data_files[9970] = "test_data_9970.txt";
test_data_files[9971] = "test_data_9971.txt";
test_data_files[9972] = "test_data_9972.txt";
test_data_files[9973] = "test_data_9973.txt";
test_data_files[9974] = "test_data_9974.txt";
test_data_files[9975] = "test_data_9975.txt";
test_data_files[9976] = "test_data_9976.txt";
test_data_files[9977] = "test_data_9977.txt";
test_data_files[9978] = "test_data_9978.txt";
test_data_files[9979] = "test_data_9979.txt";
test_data_files[9980] = "test_data_9980.txt";
test_data_files[9981] = "test_data_9981.txt";
test_data_files[9982] = "test_data_9982.txt";
test_data_files[9983] = "test_data_9983.txt";
test_data_files[9984] = "test_data_9984.txt";
test_data_files[9985] = "test_data_9985.txt";
test_data_files[9986] = "test_data_9986.txt";
test_data_files[9987] = "test_data_9987.txt";
test_data_files[9988] = "test_data_9988.txt";
test_data_files[9989] = "test_data_9989.txt";
test_data_files[9990] = "test_data_9990.txt";
test_data_files[9991] = "test_data_9991.txt";
test_data_files[9992] = "test_data_9992.txt";
test_data_files[9993] = "test_data_9993.txt";
test_data_files[9994] = "test_data_9994.txt";
test_data_files[9995] = "test_data_9995.txt";
test_data_files[9996] = "test_data_9996.txt";
test_data_files[9997] = "test_data_9997.txt";
test_data_files[9998] = "test_data_9998.txt";

    end
    
    task sendData(input [8*20-1:0] file_name);
    integer t;
    begin
        $readmemb(file_name, in_mem);
        @(posedge clock);
        @(posedge clock);
        @(posedge clock);
        for (t=0; t<784; t=t+1) begin
            @(posedge clock);
            in <= in_mem[t];
            in_valid <= 1;
        end 
        @(posedge clock);
        in_valid <= 0;
        expected = in_mem[t];
    end
    endtask
   
    integer testDataCount;
    integer start;
    initial
    begin
        reset = 0;
        in_valid = 0;
        #100;
        reset = 1;
        #100
        writeAxi(28,0); // Clear soft reset
        start = $time;
        `ifndef pretrained
            configWeights();
            configBias();
        `endif
        $display("Configuration completed",,,,$time-start,,"ns");
        start = $time;
        for(testDataCount=0; testDataCount<`MaxTestSamples; testDataCount=testDataCount+1)
        begin
            sendData(test_data_files[testDataCount]);
            @(posedge intr);
            readAxi(8);
            if(axiRdData==expected)
                right = right+1;
            $display("%0d. Accuracy: %f, Detected number: %0x, Expected: %x", testDataCount+1, right*100.0/(testDataCount+1), axiRdData, expected);
        end
        $display("Accuracy: %f", right*100.0/testDataCount);
        $stop;
    end
endmodule